magic
tech gf180mcuC
magscale 1 5
timestamp 1665299795
<< error_s >>
rect -5062 3782 -4598 3802
rect -5062 3774 -5042 3782
rect -5034 3774 -5006 3782
rect -4958 3774 -4930 3782
rect -4882 3774 -4854 3782
rect -4806 3774 -4778 3782
rect -4730 3774 -4702 3782
rect -4654 3774 -4626 3782
rect -4618 3774 -4598 3782
rect -5034 3746 -4986 3774
rect -4958 3746 -4910 3774
rect -4882 3746 -4834 3774
rect -4806 3746 -4758 3774
rect -4730 3746 -4682 3774
rect -4654 3746 -4598 3774
rect -5062 3698 -5042 3726
rect -5034 3698 -5006 3718
rect -4958 3698 -4930 3718
rect -4882 3698 -4854 3718
rect -4806 3698 -4778 3718
rect -4730 3698 -4702 3718
rect -4654 3698 -4626 3718
rect -4618 3698 -4598 3726
rect -5034 3670 -4986 3698
rect -4958 3670 -4910 3698
rect -4882 3670 -4834 3698
rect -4806 3670 -4758 3698
rect -4730 3670 -4682 3698
rect -4654 3670 -4598 3698
rect -5062 3622 -5042 3650
rect -5034 3622 -5006 3642
rect -4958 3622 -4930 3642
rect -4882 3622 -4854 3642
rect -4806 3622 -4778 3642
rect -4730 3622 -4702 3642
rect -4654 3622 -4626 3642
rect -4618 3622 -4598 3650
rect -5034 3594 -4986 3622
rect -4958 3594 -4910 3622
rect -4882 3594 -4834 3622
rect -4806 3594 -4758 3622
rect -4730 3594 -4682 3622
rect -4654 3594 -4598 3622
rect -5062 3546 -5042 3574
rect -5034 3546 -5006 3566
rect -4958 3546 -4930 3566
rect -4882 3546 -4854 3566
rect -4806 3546 -4778 3566
rect -4730 3546 -4702 3566
rect -4654 3546 -4626 3566
rect -4618 3546 -4598 3574
rect -5034 3518 -4986 3546
rect -4958 3518 -4910 3546
rect -4882 3518 -4834 3546
rect -4806 3518 -4758 3546
rect -4730 3518 -4682 3546
rect -4654 3518 -4598 3546
rect -5062 3470 -5042 3498
rect -5034 3470 -5006 3490
rect -4958 3470 -4930 3490
rect -4882 3470 -4854 3490
rect -4806 3470 -4778 3490
rect -4730 3470 -4702 3490
rect -4654 3470 -4626 3490
rect -4618 3470 -4598 3498
rect -5034 3442 -4986 3470
rect -4958 3442 -4910 3470
rect -4882 3442 -4834 3470
rect -4806 3442 -4758 3470
rect -4730 3442 -4682 3470
rect -4654 3442 -4598 3470
rect -5062 3394 -5042 3422
rect -5034 3394 -5006 3414
rect -4958 3394 -4930 3414
rect -4882 3394 -4854 3414
rect -4806 3394 -4778 3414
rect -4730 3394 -4702 3414
rect -4654 3394 -4626 3414
rect -4618 3394 -4598 3422
rect -5034 3366 -4986 3394
rect -4958 3366 -4910 3394
rect -4882 3366 -4834 3394
rect -4806 3366 -4758 3394
rect -4730 3366 -4682 3394
rect -4654 3366 -4598 3394
rect -5062 -1258 -4598 -1238
rect -5062 -1266 -5042 -1258
rect -5034 -1266 -5006 -1258
rect -4958 -1266 -4930 -1258
rect -4882 -1266 -4854 -1258
rect -4806 -1266 -4778 -1258
rect -4730 -1266 -4702 -1258
rect -4654 -1266 -4626 -1258
rect -4618 -1266 -4598 -1258
rect -5034 -1294 -4986 -1266
rect -4958 -1294 -4910 -1266
rect -4882 -1294 -4834 -1266
rect -4806 -1294 -4758 -1266
rect -4730 -1294 -4682 -1266
rect -4654 -1294 -4598 -1266
rect -5062 -1342 -5042 -1314
rect -5034 -1342 -5006 -1322
rect -4958 -1342 -4930 -1322
rect -4882 -1342 -4854 -1322
rect -4806 -1342 -4778 -1322
rect -4730 -1342 -4702 -1322
rect -4654 -1342 -4626 -1322
rect -4618 -1342 -4598 -1314
rect -5034 -1370 -4986 -1342
rect -4958 -1370 -4910 -1342
rect -4882 -1370 -4834 -1342
rect -4806 -1370 -4758 -1342
rect -4730 -1370 -4682 -1342
rect -4654 -1370 -4598 -1342
rect -5062 -1418 -5042 -1390
rect -5034 -1418 -5006 -1398
rect -4958 -1418 -4930 -1398
rect -4882 -1418 -4854 -1398
rect -4806 -1418 -4778 -1398
rect -4730 -1418 -4702 -1398
rect -4654 -1418 -4626 -1398
rect -4618 -1418 -4598 -1390
rect -5034 -1446 -4986 -1418
rect -4958 -1446 -4910 -1418
rect -4882 -1446 -4834 -1418
rect -4806 -1446 -4758 -1418
rect -4730 -1446 -4682 -1418
rect -4654 -1446 -4598 -1418
rect -5062 -1494 -5042 -1466
rect -5034 -1494 -5006 -1474
rect -4958 -1494 -4930 -1474
rect -4882 -1494 -4854 -1474
rect -4806 -1494 -4778 -1474
rect -4730 -1494 -4702 -1474
rect -4654 -1494 -4626 -1474
rect -4618 -1494 -4598 -1466
rect -5034 -1522 -4986 -1494
rect -4958 -1522 -4910 -1494
rect -4882 -1522 -4834 -1494
rect -4806 -1522 -4758 -1494
rect -4730 -1522 -4682 -1494
rect -4654 -1522 -4598 -1494
rect -5062 -1570 -5042 -1542
rect -5034 -1570 -5006 -1550
rect -4958 -1570 -4930 -1550
rect -4882 -1570 -4854 -1550
rect -4806 -1570 -4778 -1550
rect -4730 -1570 -4702 -1550
rect -4654 -1570 -4626 -1550
rect -4618 -1570 -4598 -1542
rect -5034 -1598 -4986 -1570
rect -4958 -1598 -4910 -1570
rect -4882 -1598 -4834 -1570
rect -4806 -1598 -4758 -1570
rect -4730 -1598 -4682 -1570
rect -4654 -1598 -4598 -1570
rect -5062 -1646 -5042 -1618
rect -5034 -1646 -5006 -1626
rect -4958 -1646 -4930 -1626
rect -4882 -1646 -4854 -1626
rect -4806 -1646 -4778 -1626
rect -4730 -1646 -4702 -1626
rect -4654 -1646 -4626 -1626
rect -4618 -1646 -4598 -1618
rect -5034 -1674 -4986 -1646
rect -4958 -1674 -4910 -1646
rect -4882 -1674 -4834 -1646
rect -4806 -1674 -4758 -1646
rect -4730 -1674 -4682 -1646
rect -4654 -1674 -4598 -1646
<< metal2 >>
rect -2040 1240 -1980 1260
rect -2040 1160 -2024 1240
rect -1996 1160 -1980 1240
rect -2040 1140 -1980 1160
rect -240 1240 -180 1260
rect -240 1160 -224 1240
rect -196 1160 -180 1240
rect -240 1140 -180 1160
rect 960 1240 1020 1260
rect 960 1160 976 1240
rect 1004 1160 1020 1240
rect 960 1140 1020 1160
rect 1560 1240 1620 1260
rect 1560 1160 1576 1240
rect 1604 1160 1620 1240
rect 1560 1140 1620 1160
rect 2760 1240 2820 1260
rect 2760 1160 2776 1240
rect 2804 1160 2820 1240
rect 2760 1140 2820 1160
rect 4560 1240 4620 1260
rect 4560 1160 4576 1240
rect 4604 1160 4620 1240
rect 4560 1140 4620 1160
rect 5160 1240 5220 1260
rect 5160 1160 5176 1240
rect 5204 1160 5220 1240
rect 5160 1140 5220 1160
rect 6960 1240 7020 1260
rect 6960 1160 6976 1240
rect 7004 1160 7020 1240
rect 6960 1140 7020 1160
rect 8160 1240 8220 1260
rect 8160 1160 8176 1240
rect 8204 1160 8220 1240
rect 8160 1140 8220 1160
rect 8760 1240 8820 1260
rect 8760 1160 8776 1240
rect 8804 1160 8820 1240
rect 8760 1140 8820 1160
rect 9960 1240 10020 1260
rect 9960 1160 9976 1240
rect 10004 1160 10020 1240
rect 9960 1140 10020 1160
rect 11760 1240 11820 1260
rect 11760 1160 11776 1240
rect 11804 1160 11820 1240
rect 11760 1140 11820 1160
rect -3240 1064 -3180 1080
rect -3240 1036 -3224 1064
rect -3196 1036 -3180 1064
rect -3240 1020 -3180 1036
rect -2640 1064 -2580 1080
rect -2640 1036 -2624 1064
rect -2596 1036 -2580 1064
rect -2640 1020 -2580 1036
rect 12360 1064 12420 1080
rect 12360 1036 12376 1064
rect 12404 1036 12420 1064
rect 12360 1020 12420 1036
rect 12960 1064 13020 1080
rect 12960 1036 12976 1064
rect 13004 1036 13020 1064
rect 12960 1020 13020 1036
rect -2040 940 -1980 960
rect -2040 860 -2024 940
rect -1996 860 -1980 940
rect -2040 840 -1980 860
rect -240 940 -180 960
rect -240 860 -224 940
rect -196 860 -180 940
rect -240 840 -180 860
rect 960 940 1020 960
rect 960 860 976 940
rect 1004 860 1020 940
rect 960 840 1020 860
rect 1560 940 1620 960
rect 1560 860 1576 940
rect 1604 860 1620 940
rect 1560 840 1620 860
rect 2760 940 2820 960
rect 2760 860 2776 940
rect 2804 860 2820 940
rect 2760 840 2820 860
rect 4560 940 4620 960
rect 4560 860 4576 940
rect 4604 860 4620 940
rect 4560 840 4620 860
rect 5160 940 5220 960
rect 5160 860 5176 940
rect 5204 860 5220 940
rect 5160 840 5220 860
rect 6960 940 7020 960
rect 6960 860 6976 940
rect 7004 860 7020 940
rect 6960 840 7020 860
rect 8160 940 8220 960
rect 8160 860 8176 940
rect 8204 860 8220 940
rect 8160 840 8220 860
rect 8760 940 8820 960
rect 8760 860 8776 940
rect 8804 860 8820 940
rect 8760 840 8820 860
rect 9960 940 10020 960
rect 9960 860 9976 940
rect 10004 860 10020 940
rect 9960 840 10020 860
rect 11760 940 11820 960
rect 11760 860 11776 940
rect 11804 860 11820 940
rect 11760 840 11820 860
rect -1440 160 -1380 180
rect -1440 80 -1424 160
rect -1396 80 -1380 160
rect -1440 60 -1380 80
rect -840 160 -780 180
rect -840 80 -824 160
rect -796 80 -780 160
rect -840 60 -780 80
rect 360 160 420 180
rect 360 80 376 160
rect 404 80 420 160
rect 360 60 420 80
rect 2160 160 2220 180
rect 2160 80 2176 160
rect 2204 80 2220 160
rect 2160 60 2220 80
rect 3360 160 3420 180
rect 3360 80 3376 160
rect 3404 80 3420 160
rect 3360 60 3420 80
rect 3960 160 4020 180
rect 3960 80 3976 160
rect 4004 80 4020 160
rect 3960 60 4020 80
rect 5760 160 5820 180
rect 5760 80 5776 160
rect 5804 80 5820 160
rect 5760 60 5820 80
rect 6360 160 6420 180
rect 6360 80 6376 160
rect 6404 80 6420 160
rect 6360 60 6420 80
rect 7560 160 7620 180
rect 7560 80 7576 160
rect 7604 80 7620 160
rect 7560 60 7620 80
rect 9360 160 9420 180
rect 9360 80 9376 160
rect 9404 80 9420 160
rect 9360 60 9420 80
rect 10560 160 10620 180
rect 10560 80 10576 160
rect 10604 80 10620 160
rect 10560 60 10620 80
rect 11160 160 11220 180
rect 11160 80 11176 160
rect 11204 80 11220 160
rect 11160 60 11220 80
rect -4440 -16 -4380 0
rect -4440 -44 -4424 -16
rect -4396 -44 -4380 -16
rect -4440 -60 -4380 -44
rect -3840 -16 -3780 0
rect -3840 -44 -3824 -16
rect -3796 -44 -3780 -16
rect -3840 -60 -3780 -44
rect 13560 -16 13620 0
rect 13560 -44 13576 -16
rect 13604 -44 13620 -16
rect 13560 -60 13620 -44
rect 14160 -16 14220 0
rect 14160 -44 14176 -16
rect 14204 -44 14220 -16
rect 14160 -60 14220 -44
rect -1440 -140 -1380 -120
rect -1440 -220 -1424 -140
rect -1396 -220 -1380 -140
rect -1440 -240 -1380 -220
rect -840 -140 -780 -120
rect -840 -220 -824 -140
rect -796 -220 -780 -140
rect -840 -240 -780 -220
rect 360 -140 420 -120
rect 360 -220 376 -140
rect 404 -220 420 -140
rect 360 -240 420 -220
rect 2160 -140 2220 -120
rect 2160 -220 2176 -140
rect 2204 -220 2220 -140
rect 2160 -240 2220 -220
rect 3360 -140 3420 -120
rect 3360 -220 3376 -140
rect 3404 -220 3420 -140
rect 3360 -240 3420 -220
rect 3960 -140 4020 -120
rect 3960 -220 3976 -140
rect 4004 -220 4020 -140
rect 3960 -240 4020 -220
rect 5760 -140 5820 -120
rect 5760 -220 5776 -140
rect 5804 -220 5820 -140
rect 5760 -240 5820 -220
rect 6360 -140 6420 -120
rect 6360 -220 6376 -140
rect 6404 -220 6420 -140
rect 6360 -240 6420 -220
rect 7560 -140 7620 -120
rect 7560 -220 7576 -140
rect 7604 -220 7620 -140
rect 7560 -240 7620 -220
rect 9360 -140 9420 -120
rect 9360 -220 9376 -140
rect 9404 -220 9420 -140
rect 9360 -240 9420 -220
rect 10560 -140 10620 -120
rect 10560 -220 10576 -140
rect 10604 -220 10620 -140
rect 10560 -240 10620 -220
rect 11160 -140 11220 -120
rect 11160 -220 11176 -140
rect 11204 -220 11220 -140
rect 11160 -240 11220 -220
<< via2 >>
rect -2024 1160 -1996 1240
rect -224 1160 -196 1240
rect 976 1160 1004 1240
rect 1576 1160 1604 1240
rect 2776 1160 2804 1240
rect 4576 1160 4604 1240
rect 5176 1160 5204 1240
rect 6976 1160 7004 1240
rect 8176 1160 8204 1240
rect 8776 1160 8804 1240
rect 9976 1160 10004 1240
rect 11776 1160 11804 1240
rect -3224 1036 -3196 1064
rect -2624 1036 -2596 1064
rect 12376 1036 12404 1064
rect 12976 1036 13004 1064
rect -2024 860 -1996 940
rect -224 860 -196 940
rect 976 860 1004 940
rect 1576 860 1604 940
rect 2776 860 2804 940
rect 4576 860 4604 940
rect 5176 860 5204 940
rect 6976 860 7004 940
rect 8176 860 8204 940
rect 8776 860 8804 940
rect 9976 860 10004 940
rect 11776 860 11804 940
rect -1424 80 -1396 160
rect -824 80 -796 160
rect 376 80 404 160
rect 2176 80 2204 160
rect 3376 80 3404 160
rect 3976 80 4004 160
rect 5776 80 5804 160
rect 6376 80 6404 160
rect 7576 80 7604 160
rect 9376 80 9404 160
rect 10576 80 10604 160
rect 11176 80 11204 160
rect -4424 -44 -4396 -16
rect -3824 -44 -3796 -16
rect 13576 -44 13604 -16
rect 14176 -44 14204 -16
rect -1424 -220 -1396 -140
rect -824 -220 -796 -140
rect 376 -220 404 -140
rect 2176 -220 2204 -140
rect 3376 -220 3404 -140
rect 3976 -220 4004 -140
rect 5776 -220 5804 -140
rect 6376 -220 6404 -140
rect 7576 -220 7604 -140
rect 9376 -220 9404 -140
rect 10576 -220 10604 -140
rect 11176 -220 11204 -140
<< mimcap >>
rect -5100 3782 14880 4020
rect -5100 3358 -5042 3782
rect -4618 3358 14880 3782
rect -5100 3300 14880 3358
rect -5100 -1258 14880 -1200
rect -5100 -1682 -5042 -1258
rect -4618 -1682 14880 -1258
rect -5100 -1920 14880 -1682
<< mimcapcontact >>
rect -5042 3358 -4618 3782
rect -5042 -1682 -4618 -1258
<< metal3 >>
rect -5220 2460 -5160 2760
rect -5220 2190 -5160 2280
rect -5220 2100 -5160 2160
rect -5220 1440 -5160 1500
rect -5520 1225 -5160 1260
rect -5520 1145 -5504 1225
rect -5476 1145 -5264 1225
rect -5236 1145 -5160 1225
rect -5520 1110 -5160 1145
rect -2040 1240 -1980 1260
rect -2040 1160 -2024 1240
rect -1996 1160 -1980 1240
rect -2040 1140 -1980 1160
rect -720 1240 -660 1260
rect -720 1160 -704 1240
rect -676 1160 -660 1240
rect -720 1140 -660 1160
rect -360 1240 -300 1260
rect -360 1160 -344 1240
rect -316 1160 -300 1240
rect -360 1140 -300 1160
rect -240 1240 -180 1260
rect -240 1160 -224 1240
rect -196 1160 -180 1240
rect -240 1140 -180 1160
rect 960 1240 1020 1260
rect 960 1160 976 1240
rect 1004 1160 1020 1240
rect 960 1140 1020 1160
rect 1560 1240 1620 1260
rect 1560 1160 1576 1240
rect 1604 1160 1620 1240
rect 1560 1140 1620 1160
rect 2760 1240 2820 1260
rect 2760 1160 2776 1240
rect 2804 1160 2820 1240
rect 2760 1140 2820 1160
rect 2880 1240 2940 1260
rect 2880 1160 2896 1240
rect 2924 1160 2940 1240
rect 2880 1140 2940 1160
rect 3240 1240 3300 1260
rect 3240 1160 3256 1240
rect 3284 1160 3300 1240
rect 3240 1140 3300 1160
rect 4560 1240 4620 1260
rect 4560 1160 4576 1240
rect 4604 1160 4620 1240
rect 4560 1140 4620 1160
rect 5160 1240 5220 1260
rect 5160 1160 5176 1240
rect 5204 1160 5220 1240
rect 5160 1140 5220 1160
rect 6480 1240 6540 1260
rect 6480 1160 6496 1240
rect 6524 1160 6540 1240
rect 6480 1140 6540 1160
rect 6840 1240 6900 1260
rect 6840 1160 6856 1240
rect 6884 1160 6900 1240
rect 6840 1140 6900 1160
rect 6960 1240 7020 1260
rect 6960 1160 6976 1240
rect 7004 1160 7020 1240
rect 6960 1140 7020 1160
rect 8160 1240 8220 1260
rect 8160 1160 8176 1240
rect 8204 1160 8220 1240
rect 8160 1140 8220 1160
rect 8760 1240 8820 1260
rect 8760 1160 8776 1240
rect 8804 1160 8820 1240
rect 8760 1140 8820 1160
rect 9960 1240 10020 1260
rect 9960 1160 9976 1240
rect 10004 1160 10020 1240
rect 9960 1140 10020 1160
rect 10080 1240 10140 1260
rect 10080 1160 10096 1240
rect 10124 1160 10140 1240
rect 10080 1140 10140 1160
rect 10440 1240 10500 1260
rect 10440 1160 10456 1240
rect 10484 1160 10500 1240
rect 10440 1140 10500 1160
rect 11760 1240 11820 1260
rect 11760 1160 11776 1240
rect 11804 1160 11820 1240
rect 11760 1140 11820 1160
rect -5520 1064 -5160 1080
rect -5520 1036 -5384 1064
rect -5356 1036 -5160 1064
rect -5520 1020 -5160 1036
rect -3720 1064 -3660 1080
rect -3720 1036 -3704 1064
rect -3676 1036 -3660 1064
rect -3720 1020 -3660 1036
rect -3360 1064 -3300 1080
rect -3360 1036 -3344 1064
rect -3316 1036 -3300 1064
rect -3360 1020 -3300 1036
rect -3240 1064 -3180 1080
rect -3240 1036 -3224 1064
rect -3196 1036 -3180 1064
rect -3240 1020 -3180 1036
rect -2640 1064 -2580 1080
rect -2640 1036 -2624 1064
rect -2596 1036 -2580 1064
rect -2640 1020 -2580 1036
rect -2160 1064 -2100 1080
rect -2160 1036 -2144 1064
rect -2116 1036 -2100 1064
rect -2160 1020 -2100 1036
rect 1080 1064 1140 1080
rect 1080 1036 1096 1064
rect 1124 1036 1140 1064
rect 1080 1020 1140 1036
rect 1440 1064 1500 1080
rect 1440 1036 1456 1064
rect 1484 1036 1500 1064
rect 1440 1020 1500 1036
rect 4680 1064 4740 1080
rect 4680 1036 4696 1064
rect 4724 1036 4740 1064
rect 4680 1020 4740 1036
rect 5040 1064 5100 1080
rect 5040 1036 5056 1064
rect 5084 1036 5100 1064
rect 5040 1020 5100 1036
rect 8280 1064 8340 1080
rect 8280 1036 8296 1064
rect 8324 1036 8340 1064
rect 8280 1020 8340 1036
rect 8640 1064 8700 1080
rect 8640 1036 8656 1064
rect 8684 1036 8700 1064
rect 8640 1020 8700 1036
rect 11880 1064 11940 1080
rect 11880 1036 11896 1064
rect 11924 1036 11940 1064
rect 11880 1020 11940 1036
rect 12360 1064 12420 1080
rect 12360 1036 12376 1064
rect 12404 1036 12420 1064
rect 12360 1020 12420 1036
rect 12960 1064 13020 1080
rect 12960 1036 12976 1064
rect 13004 1036 13020 1064
rect 12960 1020 13020 1036
rect 13080 1064 13140 1080
rect 13080 1036 13096 1064
rect 13124 1036 13140 1064
rect 13080 1020 13140 1036
rect 13440 1064 13500 1080
rect 13440 1036 13456 1064
rect 13484 1036 13500 1064
rect 13440 1020 13500 1036
rect -5520 955 -5160 990
rect -5520 875 -5504 955
rect -5476 875 -5264 955
rect -5236 875 -5160 955
rect -5520 840 -5160 875
rect -2040 940 -1980 960
rect -2040 860 -2024 940
rect -1996 860 -1980 940
rect -2040 840 -1980 860
rect -720 940 -660 960
rect -720 860 -704 940
rect -676 860 -660 940
rect -720 840 -660 860
rect -360 940 -300 960
rect -360 860 -344 940
rect -316 860 -300 940
rect -360 840 -300 860
rect -240 940 -180 960
rect -240 860 -224 940
rect -196 860 -180 940
rect -240 840 -180 860
rect 960 940 1020 960
rect 960 860 976 940
rect 1004 860 1020 940
rect 960 840 1020 860
rect 1560 940 1620 960
rect 1560 860 1576 940
rect 1604 860 1620 940
rect 1560 840 1620 860
rect 2760 940 2820 960
rect 2760 860 2776 940
rect 2804 860 2820 940
rect 2760 840 2820 860
rect 2880 940 2940 960
rect 2880 860 2896 940
rect 2924 860 2940 940
rect 2880 840 2940 860
rect 3240 940 3300 960
rect 3240 860 3256 940
rect 3284 860 3300 940
rect 3240 840 3300 860
rect 4560 940 4620 960
rect 4560 860 4576 940
rect 4604 860 4620 940
rect 4560 840 4620 860
rect 5160 940 5220 960
rect 5160 860 5176 940
rect 5204 860 5220 940
rect 5160 840 5220 860
rect 6480 940 6540 960
rect 6480 860 6496 940
rect 6524 860 6540 940
rect 6480 840 6540 860
rect 6840 940 6900 960
rect 6840 860 6856 940
rect 6884 860 6900 940
rect 6840 840 6900 860
rect 6960 940 7020 960
rect 6960 860 6976 940
rect 7004 860 7020 940
rect 6960 840 7020 860
rect 8160 940 8220 960
rect 8160 860 8176 940
rect 8204 860 8220 940
rect 8160 840 8220 860
rect 8760 940 8820 960
rect 8760 860 8776 940
rect 8804 860 8820 940
rect 8760 840 8820 860
rect 9960 940 10020 960
rect 9960 860 9976 940
rect 10004 860 10020 940
rect 9960 840 10020 860
rect 10080 940 10140 960
rect 10080 860 10096 940
rect 10124 860 10140 940
rect 10080 840 10140 860
rect 10440 940 10500 960
rect 10440 860 10456 940
rect 10484 860 10500 940
rect 10440 840 10500 860
rect 11760 940 11820 960
rect 11760 860 11776 940
rect 11804 860 11820 940
rect 11760 840 11820 860
rect -5220 600 -5160 660
rect -4560 644 -4500 660
rect -4560 616 -4544 644
rect -4516 616 -4500 644
rect -4560 600 -4500 616
rect -4320 644 -4260 660
rect -4320 616 -4304 644
rect -4276 616 -4260 644
rect -4320 600 -4260 616
rect -1920 644 -1860 660
rect -1920 616 -1904 644
rect -1876 616 -1860 644
rect -1920 600 -1860 616
rect 840 644 900 660
rect 840 616 856 644
rect 884 616 900 644
rect 840 600 900 616
rect 1680 644 1740 660
rect 1680 616 1696 644
rect 1724 616 1740 644
rect 1680 600 1740 616
rect 4440 644 4500 660
rect 4440 616 4456 644
rect 4484 616 4500 644
rect 4440 600 4500 616
rect 5280 644 5340 660
rect 5280 616 5296 644
rect 5324 616 5340 644
rect 5280 600 5340 616
rect 8040 644 8100 660
rect 8040 616 8056 644
rect 8084 616 8100 644
rect 8040 600 8100 616
rect 8880 644 8940 660
rect 8880 616 8896 644
rect 8924 616 8940 644
rect 8880 600 8940 616
rect 11640 644 11700 660
rect 11640 616 11656 644
rect 11684 616 11700 644
rect 11640 600 11700 616
rect 14040 644 14100 660
rect 14040 616 14056 644
rect 14084 616 14100 644
rect 14040 600 14100 616
rect 14280 644 14340 660
rect 14280 616 14296 644
rect 14324 616 14340 644
rect 14280 600 14340 616
rect -5220 360 -5160 420
rect -2760 404 -2700 420
rect -2760 376 -2744 404
rect -2716 376 -2700 404
rect -2760 360 -2700 376
rect -2520 404 -2460 420
rect -2520 376 -2504 404
rect -2476 376 -2460 404
rect -2520 360 -2460 376
rect -1560 404 -1500 420
rect -1560 376 -1544 404
rect -1516 376 -1500 404
rect -1560 360 -1500 376
rect 480 404 540 420
rect 480 376 496 404
rect 524 376 540 404
rect 480 360 540 376
rect 2040 404 2100 420
rect 2040 376 2056 404
rect 2084 376 2100 404
rect 2040 360 2100 376
rect 4080 404 4140 420
rect 4080 376 4096 404
rect 4124 376 4140 404
rect 4080 360 4140 376
rect 5640 404 5700 420
rect 5640 376 5656 404
rect 5684 376 5700 404
rect 5640 360 5700 376
rect 7680 404 7740 420
rect 7680 376 7696 404
rect 7724 376 7740 404
rect 7680 360 7740 376
rect 9240 404 9300 420
rect 9240 376 9256 404
rect 9284 376 9300 404
rect 9240 360 9300 376
rect 11280 404 11340 420
rect 11280 376 11296 404
rect 11324 376 11340 404
rect 11280 360 11340 376
rect 12240 404 12300 420
rect 12240 376 12256 404
rect 12284 376 12300 404
rect 12240 360 12300 376
rect 12480 404 12540 420
rect 12480 376 12496 404
rect 12524 376 12540 404
rect 12480 360 12540 376
rect -5520 145 -5160 180
rect -5520 65 -5504 145
rect -5476 65 -5264 145
rect -5236 65 -5160 145
rect -5520 30 -5160 65
rect -1440 160 -1380 180
rect -1440 80 -1424 160
rect -1396 80 -1380 160
rect -1440 60 -1380 80
rect -960 160 -900 180
rect -960 80 -944 160
rect -916 80 -900 160
rect -960 60 -900 80
rect -840 160 -780 180
rect -840 80 -824 160
rect -796 80 -780 160
rect -840 60 -780 80
rect -120 160 -60 180
rect -120 80 -104 160
rect -76 80 -60 160
rect -120 60 -60 80
rect 360 160 420 180
rect 360 80 376 160
rect 404 80 420 160
rect 360 60 420 80
rect 2160 160 2220 180
rect 2160 80 2176 160
rect 2204 80 2220 160
rect 2160 60 2220 80
rect 2640 160 2700 180
rect 2640 80 2656 160
rect 2684 80 2700 160
rect 2640 60 2700 80
rect 3360 160 3420 180
rect 3360 80 3376 160
rect 3404 80 3420 160
rect 3360 60 3420 80
rect 3480 160 3540 180
rect 3480 80 3496 160
rect 3524 80 3540 160
rect 3480 60 3540 80
rect 3960 160 4020 180
rect 3960 80 3976 160
rect 4004 80 4020 160
rect 3960 60 4020 80
rect 5760 160 5820 180
rect 5760 80 5776 160
rect 5804 80 5820 160
rect 5760 60 5820 80
rect 6240 160 6300 180
rect 6240 80 6256 160
rect 6284 80 6300 160
rect 6240 60 6300 80
rect 6360 160 6420 180
rect 6360 80 6376 160
rect 6404 80 6420 160
rect 6360 60 6420 80
rect 7080 160 7140 180
rect 7080 80 7096 160
rect 7124 80 7140 160
rect 7080 60 7140 80
rect 7560 160 7620 180
rect 7560 80 7576 160
rect 7604 80 7620 160
rect 7560 60 7620 80
rect 9360 160 9420 180
rect 9360 80 9376 160
rect 9404 80 9420 160
rect 9360 60 9420 80
rect 9840 160 9900 180
rect 9840 80 9856 160
rect 9884 80 9900 160
rect 9840 60 9900 80
rect 10560 160 10620 180
rect 10560 80 10576 160
rect 10604 80 10620 160
rect 10560 60 10620 80
rect 10680 160 10740 180
rect 10680 80 10696 160
rect 10724 80 10740 160
rect 10680 60 10740 80
rect 11160 160 11220 180
rect 11160 80 11176 160
rect 11204 80 11220 160
rect 11160 60 11220 80
rect -5520 -16 -5160 0
rect -5520 -44 -5384 -16
rect -5356 -44 -5160 -16
rect -5520 -60 -5160 -44
rect -4440 -16 -4380 0
rect -4440 -44 -4424 -16
rect -4396 -44 -4380 -16
rect -4440 -60 -4380 -44
rect -3960 -16 -3900 0
rect -3960 -44 -3944 -16
rect -3916 -44 -3900 -16
rect -3960 -60 -3900 -44
rect -3840 -16 -3780 0
rect -3840 -44 -3824 -16
rect -3796 -44 -3780 -16
rect -3840 -60 -3780 -44
rect -3120 -16 -3060 0
rect -3120 -44 -3104 -16
rect -3076 -44 -3060 -16
rect -3120 -60 -3060 -44
rect -1320 -16 -1260 0
rect -1320 -44 -1304 -16
rect -1276 -44 -1260 -16
rect -1320 -60 -1260 -44
rect 240 -16 300 0
rect 240 -44 256 -16
rect 284 -44 300 -16
rect 240 -60 300 -44
rect 2280 -16 2340 0
rect 2280 -44 2296 -16
rect 2324 -44 2340 -16
rect 2280 -60 2340 -44
rect 3840 -16 3900 0
rect 3840 -44 3856 -16
rect 3884 -44 3900 -16
rect 3840 -60 3900 -44
rect 5880 -16 5940 0
rect 5880 -44 5896 -16
rect 5924 -44 5940 -16
rect 5880 -60 5940 -44
rect 7440 -16 7500 0
rect 7440 -44 7456 -16
rect 7484 -44 7500 -16
rect 7440 -60 7500 -44
rect 9480 -16 9540 0
rect 9480 -44 9496 -16
rect 9524 -44 9540 -16
rect 9480 -60 9540 -44
rect 11040 -16 11100 0
rect 11040 -44 11056 -16
rect 11084 -44 11100 -16
rect 11040 -60 11100 -44
rect 12840 -16 12900 0
rect 12840 -44 12856 -16
rect 12884 -44 12900 -16
rect 12840 -60 12900 -44
rect 13560 -16 13620 0
rect 13560 -44 13576 -16
rect 13604 -44 13620 -16
rect 13560 -60 13620 -44
rect 13680 -16 13740 0
rect 13680 -44 13696 -16
rect 13724 -44 13740 -16
rect 13680 -60 13740 -44
rect 14160 -16 14220 0
rect 14160 -44 14176 -16
rect 14204 -44 14220 -16
rect 14160 -60 14220 -44
rect -5520 -125 -5160 -90
rect -5520 -205 -5504 -125
rect -5476 -205 -5264 -125
rect -5236 -205 -5160 -125
rect -5520 -240 -5160 -205
rect -1440 -140 -1380 -120
rect -1440 -220 -1424 -140
rect -1396 -220 -1380 -140
rect -1440 -240 -1380 -220
rect -960 -140 -900 -120
rect -960 -220 -944 -140
rect -916 -220 -900 -140
rect -960 -240 -900 -220
rect -840 -140 -780 -120
rect -840 -220 -824 -140
rect -796 -220 -780 -140
rect -840 -240 -780 -220
rect -120 -140 -60 -120
rect -120 -220 -104 -140
rect -76 -220 -60 -140
rect -120 -240 -60 -220
rect 360 -140 420 -120
rect 360 -220 376 -140
rect 404 -220 420 -140
rect 360 -240 420 -220
rect 2160 -140 2220 -120
rect 2160 -220 2176 -140
rect 2204 -220 2220 -140
rect 2160 -240 2220 -220
rect 2640 -140 2700 -120
rect 2640 -220 2656 -140
rect 2684 -220 2700 -140
rect 2640 -240 2700 -220
rect 3360 -140 3420 -120
rect 3360 -220 3376 -140
rect 3404 -220 3420 -140
rect 3360 -240 3420 -220
rect 3480 -140 3540 -120
rect 3480 -220 3496 -140
rect 3524 -220 3540 -140
rect 3480 -240 3540 -220
rect 3960 -140 4020 -120
rect 3960 -220 3976 -140
rect 4004 -220 4020 -140
rect 3960 -240 4020 -220
rect 5760 -140 5820 -120
rect 5760 -220 5776 -140
rect 5804 -220 5820 -140
rect 5760 -240 5820 -220
rect 6240 -140 6300 -120
rect 6240 -220 6256 -140
rect 6284 -220 6300 -140
rect 6240 -240 6300 -220
rect 6360 -140 6420 -120
rect 6360 -220 6376 -140
rect 6404 -220 6420 -140
rect 6360 -240 6420 -220
rect 7080 -140 7140 -120
rect 7080 -220 7096 -140
rect 7124 -220 7140 -140
rect 7080 -240 7140 -220
rect 7560 -140 7620 -120
rect 7560 -220 7576 -140
rect 7604 -220 7620 -140
rect 7560 -240 7620 -220
rect 9360 -140 9420 -120
rect 9360 -220 9376 -140
rect 9404 -220 9420 -140
rect 9360 -240 9420 -220
rect 9840 -140 9900 -120
rect 9840 -220 9856 -140
rect 9884 -220 9900 -140
rect 9840 -240 9900 -220
rect 10560 -140 10620 -120
rect 10560 -220 10576 -140
rect 10604 -220 10620 -140
rect 10560 -240 10620 -220
rect 10680 -140 10740 -120
rect 10680 -220 10696 -140
rect 10724 -220 10740 -140
rect 10680 -240 10740 -220
rect 11160 -140 11220 -120
rect 11160 -220 11176 -140
rect 11204 -220 11220 -140
rect 11160 -240 11220 -220
rect -5220 -840 -5160 -540
<< via3 >>
rect -5504 1145 -5476 1225
rect -5264 1145 -5236 1225
rect -704 1160 -676 1240
rect -344 1160 -316 1240
rect 2896 1160 2924 1240
rect 3256 1160 3284 1240
rect 6496 1160 6524 1240
rect 6856 1160 6884 1240
rect 10096 1160 10124 1240
rect 10456 1160 10484 1240
rect -5384 1036 -5356 1064
rect -3704 1036 -3676 1064
rect -3344 1036 -3316 1064
rect -2144 1036 -2116 1064
rect 1096 1036 1124 1064
rect 1456 1036 1484 1064
rect 4696 1036 4724 1064
rect 5056 1036 5084 1064
rect 8296 1036 8324 1064
rect 8656 1036 8684 1064
rect 11896 1036 11924 1064
rect 13096 1036 13124 1064
rect 13456 1036 13484 1064
rect -5504 875 -5476 955
rect -5264 875 -5236 955
rect -704 860 -676 940
rect -344 860 -316 940
rect 2896 860 2924 940
rect 3256 860 3284 940
rect 6496 860 6524 940
rect 6856 860 6884 940
rect 10096 860 10124 940
rect 10456 860 10484 940
rect -4544 616 -4516 644
rect -4304 616 -4276 644
rect -1904 616 -1876 644
rect 856 616 884 644
rect 1696 616 1724 644
rect 4456 616 4484 644
rect 5296 616 5324 644
rect 8056 616 8084 644
rect 8896 616 8924 644
rect 11656 616 11684 644
rect 14056 616 14084 644
rect 14296 616 14324 644
rect -2744 376 -2716 404
rect -2504 376 -2476 404
rect -1544 376 -1516 404
rect 496 376 524 404
rect 2056 376 2084 404
rect 4096 376 4124 404
rect 5656 376 5684 404
rect 7696 376 7724 404
rect 9256 376 9284 404
rect 11296 376 11324 404
rect 12256 376 12284 404
rect 12496 376 12524 404
rect -5504 65 -5476 145
rect -5264 65 -5236 145
rect -944 80 -916 160
rect -104 80 -76 160
rect 2656 80 2684 160
rect 3496 80 3524 160
rect 6256 80 6284 160
rect 7096 80 7124 160
rect 9856 80 9884 160
rect 10696 80 10724 160
rect -5384 -44 -5356 -16
rect -3944 -44 -3916 -16
rect -3104 -44 -3076 -16
rect -1304 -44 -1276 -16
rect 256 -44 284 -16
rect 2296 -44 2324 -16
rect 3856 -44 3884 -16
rect 5896 -44 5924 -16
rect 7456 -44 7484 -16
rect 9496 -44 9524 -16
rect 11056 -44 11084 -16
rect 12856 -44 12884 -16
rect 13696 -44 13724 -16
rect -5504 -205 -5476 -125
rect -5264 -205 -5236 -125
rect -944 -220 -916 -140
rect -104 -220 -76 -140
rect 2656 -220 2684 -140
rect 3496 -220 3524 -140
rect 6256 -220 6284 -140
rect 7096 -220 7124 -140
rect 9856 -220 9884 -140
rect 10696 -220 10724 -140
<< metal4 >>
rect -5160 4020 14940 4080
rect -5520 3284 -5460 3360
rect -5520 3256 -5504 3284
rect -5476 3256 -5460 3284
rect -5520 3044 -5460 3256
rect -5520 3016 -5504 3044
rect -5476 3016 -5460 3044
rect -5520 1225 -5460 3016
rect -5520 1145 -5504 1225
rect -5476 1145 -5460 1225
rect -5520 955 -5460 1145
rect -5520 875 -5504 955
rect -5476 875 -5460 955
rect -5520 840 -5460 875
rect -5400 3164 -5340 3360
rect -5400 3136 -5384 3164
rect -5356 3136 -5340 3164
rect -5400 1064 -5340 3136
rect -5400 1036 -5384 1064
rect -5356 1036 -5340 1064
rect -5400 840 -5340 1036
rect -5280 3284 -5220 3360
rect -5280 3256 -5264 3284
rect -5236 3256 -5220 3284
rect -5280 3044 -5220 3256
rect -5160 3300 -5100 4020
rect 14880 3300 14940 4020
rect -5160 3164 14940 3300
rect -5160 3136 -5082 3164
rect 14862 3136 14940 3164
rect -5160 3120 14940 3136
rect -5280 3016 -5264 3044
rect -5236 3016 -5220 3044
rect -5280 1225 -5220 3016
rect -5280 1145 -5264 1225
rect -5236 1145 -5220 1225
rect -5280 955 -5220 1145
rect -720 1240 -660 1260
rect -720 1160 -704 1240
rect -676 1160 -660 1240
rect -720 1140 -660 1160
rect -360 1240 -300 1260
rect -360 1160 -344 1240
rect -316 1160 -300 1240
rect -360 1140 -300 1160
rect 2880 1240 2940 1260
rect 2880 1160 2896 1240
rect 2924 1160 2940 1240
rect 2880 1140 2940 1160
rect 3240 1240 3300 1260
rect 3240 1160 3256 1240
rect 3284 1160 3300 1240
rect 3240 1140 3300 1160
rect 6480 1240 6540 1260
rect 6480 1160 6496 1240
rect 6524 1160 6540 1240
rect 6480 1140 6540 1160
rect 6840 1240 6900 1260
rect 6840 1160 6856 1240
rect 6884 1160 6900 1240
rect 6840 1140 6900 1160
rect 10080 1240 10140 1260
rect 10080 1160 10096 1240
rect 10124 1160 10140 1240
rect 10080 1140 10140 1160
rect 10440 1240 10500 1260
rect 10440 1160 10456 1240
rect 10484 1160 10500 1240
rect 10440 1140 10500 1160
rect -3720 1064 -3660 1080
rect -3720 1036 -3704 1064
rect -3676 1036 -3660 1064
rect -3720 1020 -3660 1036
rect -3360 1064 -3300 1080
rect -3360 1036 -3344 1064
rect -3316 1036 -3300 1064
rect -3360 1020 -3300 1036
rect -2160 1064 -2100 1080
rect -2160 1036 -2144 1064
rect -2116 1036 -2100 1064
rect -2160 1020 -2100 1036
rect 1080 1064 1140 1080
rect 1080 1036 1096 1064
rect 1124 1036 1140 1064
rect 1080 1020 1140 1036
rect 1440 1064 1500 1080
rect 1440 1036 1456 1064
rect 1484 1036 1500 1064
rect 1440 1020 1500 1036
rect 4680 1064 4740 1080
rect 4680 1036 4696 1064
rect 4724 1036 4740 1064
rect 4680 1020 4740 1036
rect 5040 1064 5100 1080
rect 5040 1036 5056 1064
rect 5084 1036 5100 1064
rect 5040 1020 5100 1036
rect 8280 1064 8340 1080
rect 8280 1036 8296 1064
rect 8324 1036 8340 1064
rect 8280 1020 8340 1036
rect 8640 1064 8700 1080
rect 8640 1036 8656 1064
rect 8684 1036 8700 1064
rect 8640 1020 8700 1036
rect 11880 1064 11940 1080
rect 11880 1036 11896 1064
rect 11924 1036 11940 1064
rect 11880 1020 11940 1036
rect 13080 1064 13140 1080
rect 13080 1036 13096 1064
rect 13124 1036 13140 1064
rect 13080 1020 13140 1036
rect 13440 1064 13500 1080
rect 13440 1036 13456 1064
rect 13484 1036 13500 1064
rect 13440 1020 13500 1036
rect -5280 875 -5264 955
rect -5236 875 -5220 955
rect -5280 840 -5220 875
rect -720 940 -660 960
rect -720 860 -704 940
rect -676 860 -660 940
rect -720 840 -660 860
rect -360 940 -300 960
rect -360 860 -344 940
rect -316 860 -300 940
rect -360 840 -300 860
rect 2880 940 2940 960
rect 2880 860 2896 940
rect 2924 860 2940 940
rect 2880 840 2940 860
rect 3240 940 3300 960
rect 3240 860 3256 940
rect 3284 860 3300 940
rect 3240 840 3300 860
rect 6480 940 6540 960
rect 6480 860 6496 940
rect 6524 860 6540 940
rect 6480 840 6540 860
rect 6840 940 6900 960
rect 6840 860 6856 940
rect 6884 860 6900 940
rect 6840 840 6900 860
rect 10080 940 10140 960
rect 10080 860 10096 940
rect 10124 860 10140 940
rect 10080 840 10140 860
rect 10440 940 10500 960
rect 10440 860 10456 940
rect 10484 860 10500 940
rect 10440 840 10500 860
rect -4560 644 -4500 660
rect -4560 616 -4544 644
rect -4516 616 -4500 644
rect -4560 600 -4500 616
rect -4320 644 -4260 660
rect -4320 616 -4304 644
rect -4276 616 -4260 644
rect -4320 600 -4260 616
rect -1920 644 -1860 660
rect -1920 616 -1904 644
rect -1876 616 -1860 644
rect -1920 600 -1860 616
rect 840 644 900 660
rect 840 616 856 644
rect 884 616 900 644
rect 840 600 900 616
rect 1680 644 1740 660
rect 1680 616 1696 644
rect 1724 616 1740 644
rect 1680 600 1740 616
rect 4440 644 4500 660
rect 4440 616 4456 644
rect 4484 616 4500 644
rect 4440 600 4500 616
rect 5280 644 5340 660
rect 5280 616 5296 644
rect 5324 616 5340 644
rect 5280 600 5340 616
rect 8040 644 8100 660
rect 8040 616 8056 644
rect 8084 616 8100 644
rect 8040 600 8100 616
rect 8880 644 8940 660
rect 8880 616 8896 644
rect 8924 616 8940 644
rect 8880 600 8940 616
rect 11640 644 11700 660
rect 11640 616 11656 644
rect 11684 616 11700 644
rect 11640 600 11700 616
rect 14040 644 14100 660
rect 14040 616 14056 644
rect 14084 616 14100 644
rect 14040 600 14100 616
rect 14280 644 14340 660
rect 14280 616 14296 644
rect 14324 616 14340 644
rect 14280 600 14340 616
rect -2760 404 -2700 420
rect -2760 376 -2744 404
rect -2716 376 -2700 404
rect -2760 360 -2700 376
rect -2520 404 -2460 420
rect -2520 376 -2504 404
rect -2476 376 -2460 404
rect -2520 360 -2460 376
rect -1560 404 -1500 420
rect -1560 376 -1544 404
rect -1516 376 -1500 404
rect -1560 360 -1500 376
rect 480 404 540 420
rect 480 376 496 404
rect 524 376 540 404
rect 480 360 540 376
rect 2040 404 2100 420
rect 2040 376 2056 404
rect 2084 376 2100 404
rect 2040 360 2100 376
rect 4080 404 4140 420
rect 4080 376 4096 404
rect 4124 376 4140 404
rect 4080 360 4140 376
rect 5640 404 5700 420
rect 5640 376 5656 404
rect 5684 376 5700 404
rect 5640 360 5700 376
rect 7680 404 7740 420
rect 7680 376 7696 404
rect 7724 376 7740 404
rect 7680 360 7740 376
rect 9240 404 9300 420
rect 9240 376 9256 404
rect 9284 376 9300 404
rect 9240 360 9300 376
rect 11280 404 11340 420
rect 11280 376 11296 404
rect 11324 376 11340 404
rect 11280 360 11340 376
rect 12240 404 12300 420
rect 12240 376 12256 404
rect 12284 376 12300 404
rect 12240 360 12300 376
rect 12480 404 12540 420
rect 12480 376 12496 404
rect 12524 376 12540 404
rect 12480 360 12540 376
rect -5520 145 -5460 180
rect -5520 65 -5504 145
rect -5476 65 -5460 145
rect -5520 -125 -5460 65
rect -5520 -205 -5504 -125
rect -5476 -205 -5460 -125
rect -5520 -916 -5460 -205
rect -5520 -944 -5504 -916
rect -5476 -944 -5460 -916
rect -5520 -1156 -5460 -944
rect -5520 -1184 -5504 -1156
rect -5476 -1184 -5460 -1156
rect -5520 -1260 -5460 -1184
rect -5400 -16 -5340 180
rect -5400 -44 -5384 -16
rect -5356 -44 -5340 -16
rect -5400 -1036 -5340 -44
rect -5400 -1064 -5384 -1036
rect -5356 -1064 -5340 -1036
rect -5400 -1260 -5340 -1064
rect -5280 145 -5220 180
rect -5280 65 -5264 145
rect -5236 65 -5220 145
rect -5280 -125 -5220 65
rect -960 160 -900 180
rect -960 80 -944 160
rect -916 80 -900 160
rect -960 60 -900 80
rect -120 160 -60 180
rect -120 80 -104 160
rect -76 80 -60 160
rect -120 60 -60 80
rect 2640 160 2700 180
rect 2640 80 2656 160
rect 2684 80 2700 160
rect 2640 60 2700 80
rect 3480 160 3540 180
rect 3480 80 3496 160
rect 3524 80 3540 160
rect 3480 60 3540 80
rect 6240 160 6300 180
rect 6240 80 6256 160
rect 6284 80 6300 160
rect 6240 60 6300 80
rect 7080 160 7140 180
rect 7080 80 7096 160
rect 7124 80 7140 160
rect 7080 60 7140 80
rect 9840 160 9900 180
rect 9840 80 9856 160
rect 9884 80 9900 160
rect 9840 60 9900 80
rect 10680 160 10740 180
rect 10680 80 10696 160
rect 10724 80 10740 160
rect 10680 60 10740 80
rect -3960 -16 -3900 0
rect -3960 -44 -3944 -16
rect -3916 -44 -3900 -16
rect -3960 -60 -3900 -44
rect -3120 -16 -3060 0
rect -3120 -44 -3104 -16
rect -3076 -44 -3060 -16
rect -3120 -60 -3060 -44
rect -1320 -16 -1260 0
rect -1320 -44 -1304 -16
rect -1276 -44 -1260 -16
rect -1320 -60 -1260 -44
rect 240 -16 300 0
rect 240 -44 256 -16
rect 284 -44 300 -16
rect 240 -60 300 -44
rect 2280 -16 2340 0
rect 2280 -44 2296 -16
rect 2324 -44 2340 -16
rect 2280 -60 2340 -44
rect 3840 -16 3900 0
rect 3840 -44 3856 -16
rect 3884 -44 3900 -16
rect 3840 -60 3900 -44
rect 5880 -16 5940 0
rect 5880 -44 5896 -16
rect 5924 -44 5940 -16
rect 5880 -60 5940 -44
rect 7440 -16 7500 0
rect 7440 -44 7456 -16
rect 7484 -44 7500 -16
rect 7440 -60 7500 -44
rect 9480 -16 9540 0
rect 9480 -44 9496 -16
rect 9524 -44 9540 -16
rect 9480 -60 9540 -44
rect 11040 -16 11100 0
rect 11040 -44 11056 -16
rect 11084 -44 11100 -16
rect 11040 -60 11100 -44
rect 12840 -16 12900 0
rect 12840 -44 12856 -16
rect 12884 -44 12900 -16
rect 12840 -60 12900 -44
rect 13680 -16 13740 0
rect 13680 -44 13696 -16
rect 13724 -44 13740 -16
rect 13680 -60 13740 -44
rect -5280 -205 -5264 -125
rect -5236 -205 -5220 -125
rect -5280 -916 -5220 -205
rect -960 -140 -900 -120
rect -960 -220 -944 -140
rect -916 -220 -900 -140
rect -960 -240 -900 -220
rect -120 -140 -60 -120
rect -120 -220 -104 -140
rect -76 -220 -60 -140
rect -120 -240 -60 -220
rect 2640 -140 2700 -120
rect 2640 -220 2656 -140
rect 2684 -220 2700 -140
rect 2640 -240 2700 -220
rect 3480 -140 3540 -120
rect 3480 -220 3496 -140
rect 3524 -220 3540 -140
rect 3480 -240 3540 -220
rect 6240 -140 6300 -120
rect 6240 -220 6256 -140
rect 6284 -220 6300 -140
rect 6240 -240 6300 -220
rect 7080 -140 7140 -120
rect 7080 -220 7096 -140
rect 7124 -220 7140 -140
rect 7080 -240 7140 -220
rect 9840 -140 9900 -120
rect 9840 -220 9856 -140
rect 9884 -220 9900 -140
rect 9840 -240 9900 -220
rect 10680 -140 10740 -120
rect 10680 -220 10696 -140
rect 10724 -220 10740 -140
rect 10680 -240 10740 -220
rect -5280 -944 -5264 -916
rect -5236 -944 -5220 -916
rect -5280 -1156 -5220 -944
rect -5280 -1184 -5264 -1156
rect -5236 -1184 -5220 -1156
rect -5280 -1260 -5220 -1184
rect -5160 -1036 14940 -1020
rect -5160 -1064 -5082 -1036
rect 14862 -1064 14940 -1036
rect -5160 -1200 14940 -1064
rect -5160 -1920 -5100 -1200
rect 14880 -1920 14940 -1200
rect -5160 -1980 14940 -1920
<< via4 >>
rect -5504 3256 -5476 3284
rect -5504 3016 -5476 3044
rect -5384 3136 -5356 3164
rect -5264 3256 -5236 3284
rect -5082 3136 14862 3164
rect -5264 3016 -5236 3044
rect -5504 -944 -5476 -916
rect -5504 -1184 -5476 -1156
rect -5384 -1064 -5356 -1036
rect -5264 -944 -5236 -916
rect -5264 -1184 -5236 -1156
rect -5082 -1064 14862 -1036
<< metal5 >>
rect -5160 3782 14940 4080
rect -5160 3358 -5042 3782
rect -4618 3358 14940 3782
rect -5160 3300 14940 3358
rect -5580 3284 14940 3300
rect -5580 3256 -5504 3284
rect -5476 3256 -5264 3284
rect -5236 3256 14940 3284
rect -5580 3240 14940 3256
rect -5580 3164 14940 3180
rect -5580 3136 -5384 3164
rect -5356 3136 -5082 3164
rect 14862 3136 14940 3164
rect -5580 3120 14940 3136
rect -5580 3044 14940 3060
rect -5580 3016 -5504 3044
rect -5476 3016 -5264 3044
rect -5236 3016 14940 3044
rect -5580 3000 14940 3016
rect -5580 -916 14940 -900
rect -5580 -944 -5504 -916
rect -5476 -944 -5264 -916
rect -5236 -944 14940 -916
rect -5580 -960 14940 -944
rect -5580 -1036 14940 -1020
rect -5580 -1064 -5384 -1036
rect -5356 -1064 -5082 -1036
rect 14862 -1064 14940 -1036
rect -5580 -1080 14940 -1064
rect -5580 -1156 14940 -1140
rect -5580 -1184 -5504 -1156
rect -5476 -1184 -5264 -1156
rect -5236 -1184 14940 -1156
rect -5580 -1200 14940 -1184
rect -5160 -1258 14940 -1200
rect -5160 -1682 -5042 -1258
rect -4618 -1682 14940 -1258
rect -5160 -1980 14940 -1682
use nautanauta_cell#0  nautanauta_cell_0
timestamp 1665184495
transform -1 0 10920 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_1
timestamp 1665184495
transform -1 0 10320 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_2
timestamp 1665184495
transform -1 0 9120 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_3
timestamp 1665184495
transform -1 0 9720 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_4
timestamp 1665184495
transform -1 0 8520 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_5
timestamp 1665184495
transform -1 0 7920 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_6
timestamp 1665184495
transform -1 0 7320 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_7
timestamp 1665184495
transform -1 0 6720 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_8
timestamp 1665184495
transform -1 0 6120 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_9
timestamp 1665184495
transform -1 0 5520 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_10
timestamp 1665184495
transform 1 0 11460 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_11
timestamp 1665184495
transform 1 0 10860 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_12
timestamp 1665184495
transform 1 0 10260 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_13
timestamp 1665184495
transform 1 0 9060 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_14
timestamp 1665184495
transform 1 0 9660 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_15
timestamp 1665184495
transform 1 0 8460 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_16
timestamp 1665184495
transform -1 0 1320 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_17
timestamp 1665184495
transform -1 0 720 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_18
timestamp 1665184495
transform -1 0 120 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_19
timestamp 1665184495
transform -1 0 -480 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_20
timestamp 1665184495
transform -1 0 -1080 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_21
timestamp 1665184495
transform -1 0 -1680 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_22
timestamp 1665184495
transform 1 0 4260 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_23
timestamp 1665184495
transform 1 0 3660 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_24
timestamp 1665184495
transform 1 0 3060 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_25
timestamp 1665184495
transform 1 0 2460 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_26
timestamp 1665184495
transform 1 0 1860 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_27
timestamp 1665184495
transform 1 0 1260 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_28
timestamp 1665184495
transform 1 0 660 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_29
timestamp 1665184495
transform 1 0 60 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_30
timestamp 1665184495
transform 1 0 -540 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_cell#0  nautanauta_cell_31
timestamp 1665184495
transform 1 0 -1140 0 1 -180
box -3600 -660 -2940 3060
use nautanauta_edge#0  nautanauta_edge_0
timestamp 1665184495
transform -1 0 11160 0 1 -180
box -3780 -660 -3300 3060
use nautanauta_edge#0  nautanauta_edge_1
timestamp 1665184495
transform 1 0 -1380 0 1 -180
box -3780 -660 -3300 3060
<< labels >>
rlabel metal3 s -5190 1050 -5190 1050 4 xm
rlabel metal3 s -5190 -30 -5190 -30 4 xp
rlabel metal3 s -5220 360 -5160 420 4 ip
port 1 nsew
rlabel metal3 s -5220 600 -5160 660 4 im
port 2 nsew
rlabel metal3 s -5220 1200 -5160 1260 4 op
port 3 nsew
rlabel metal3 s -5220 -240 -5160 -180 4 om
port 4 nsew
rlabel metal3 s -5220 2460 -5160 2760 4 vdd
port 5 nsew
rlabel metal3 s -5220 2100 -5160 2160 4 gp
port 6 nsew
rlabel metal3 s -5220 1440 -5160 1500 4 bp
port 7 nsew
rlabel metal3 s -5220 2220 -5160 2280 4 vreg
port 8 nsew
rlabel metal3 s -5220 -840 -5160 -540 4 gnd
port 9 nsew
<< end >>
