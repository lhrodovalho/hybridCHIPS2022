magic
tech gf180mcuC
magscale 1 5
timestamp 1665184495
<< metal1 >>
rect -4620 1200 -4560 1260
rect -60 1200 0 1260
<< metal2 >>
rect -4440 1014 -4380 1020
rect -4440 726 -4424 1014
rect -4396 726 -4380 1014
rect -4440 720 -4380 726
rect -3840 1014 -3780 1020
rect -3840 726 -3824 1014
rect -3796 726 -3780 1014
rect -3840 720 -3780 726
rect -840 1014 -780 1020
rect -840 726 -824 1014
rect -796 726 -780 1014
rect -840 720 -780 726
rect -240 1014 -180 1020
rect -240 726 -224 1014
rect -196 726 -180 1014
rect -240 720 -180 726
rect -3240 54 -3180 60
rect -3240 -234 -3224 54
rect -3196 -234 -3180 54
rect -3240 -240 -3180 -234
rect -2640 54 -2580 60
rect -2640 -234 -2624 54
rect -2596 -234 -2580 54
rect -2640 -240 -2580 -234
rect -2040 54 -1980 60
rect -2040 -234 -2024 54
rect -1996 -234 -1980 54
rect -2040 -240 -1980 -234
rect -1440 54 -1380 60
rect -1440 -234 -1424 54
rect -1396 -234 -1380 54
rect -1440 -240 -1380 -234
<< via2 >>
rect -4424 726 -4396 1014
rect -3824 726 -3796 1014
rect -824 726 -796 1014
rect -224 726 -196 1014
rect -3224 -234 -3196 54
rect -2624 -234 -2596 54
rect -2024 -234 -1996 54
rect -1424 -234 -1396 54
<< metal3 >>
rect -5220 2220 -5160 2520
rect -5220 1950 -5160 2040
rect -5220 1860 -5160 1920
rect -5220 1200 -5160 1260
rect -4740 1200 -4430 1260
rect -190 1200 120 1260
rect -5220 720 -5160 1020
rect -4440 1014 -4380 1020
rect -4440 726 -4424 1014
rect -4396 726 -4380 1014
rect -4440 720 -4380 726
rect -4320 1014 -4260 1020
rect -4320 726 -4304 1014
rect -4276 726 -4260 1014
rect -4320 720 -4260 726
rect -3840 1014 -3780 1020
rect -3840 726 -3824 1014
rect -3796 726 -3780 1014
rect -3840 720 -3780 726
rect -3360 1014 -3300 1020
rect -3360 726 -3344 1014
rect -3316 726 -3300 1014
rect -3360 720 -3300 726
rect -1320 1014 -1260 1020
rect -1320 726 -1304 1014
rect -1276 726 -1260 1014
rect -1320 720 -1260 726
rect -840 1014 -780 1020
rect -840 726 -824 1014
rect -796 726 -780 1014
rect -840 720 -780 726
rect -360 1014 -300 1020
rect -360 726 -344 1014
rect -316 726 -300 1014
rect -360 720 -300 726
rect -240 1014 -180 1020
rect -240 726 -224 1014
rect -196 726 -180 1014
rect -240 720 -180 726
rect -5220 480 -5160 540
rect -4560 524 -4500 540
rect -4560 496 -4544 524
rect -4516 496 -4500 524
rect -4560 480 -4500 496
rect -3960 524 -3900 540
rect -3960 496 -3944 524
rect -3916 496 -3900 524
rect -3960 480 -3900 496
rect -720 524 -660 540
rect -720 496 -704 524
rect -676 496 -660 524
rect -720 480 -660 496
rect -120 524 -60 540
rect -120 496 -104 524
rect -76 496 -60 524
rect -120 480 -60 496
rect -5220 240 -5160 300
rect -3120 284 -3060 300
rect -3120 256 -3104 284
rect -3076 256 -3060 284
rect -3120 240 -3060 256
rect -2760 284 -2700 300
rect -2760 256 -2744 284
rect -2716 256 -2700 284
rect -2760 240 -2700 256
rect -1920 284 -1860 300
rect -1920 256 -1904 284
rect -1876 256 -1860 284
rect -1920 240 -1860 256
rect -1560 284 -1500 300
rect -1560 256 -1544 284
rect -1516 256 -1500 284
rect -1560 240 -1500 256
rect -5220 -240 -5160 60
rect -3720 54 -3660 60
rect -3720 -234 -3704 54
rect -3676 -234 -3660 54
rect -3720 -240 -3660 -234
rect -3240 54 -3180 60
rect -3240 -234 -3224 54
rect -3196 -234 -3180 54
rect -3240 -240 -3180 -234
rect -2640 54 -2580 60
rect -2640 -234 -2624 54
rect -2596 -234 -2580 54
rect -2640 -240 -2580 -234
rect -2520 54 -2460 60
rect -2520 -234 -2504 54
rect -2476 -234 -2460 54
rect -2520 -240 -2460 -234
rect -2160 54 -2100 60
rect -2160 -234 -2144 54
rect -2116 -234 -2100 54
rect -2160 -240 -2100 -234
rect -2040 54 -1980 60
rect -2040 -234 -2024 54
rect -1996 -234 -1980 54
rect -2040 -240 -1980 -234
rect -1440 54 -1380 60
rect -1440 -234 -1424 54
rect -1396 -234 -1380 54
rect -1440 -240 -1380 -234
rect -960 54 -900 60
rect -960 -234 -944 54
rect -916 -234 -900 54
rect -960 -240 -900 -234
rect -5220 -840 -5160 -540
<< via3 >>
rect -4304 726 -4276 1014
rect -3344 726 -3316 1014
rect -1304 726 -1276 1014
rect -344 726 -316 1014
rect -4544 496 -4516 524
rect -3944 496 -3916 524
rect -704 496 -676 524
rect -104 496 -76 524
rect -3104 256 -3076 284
rect -2744 256 -2716 284
rect -1904 256 -1876 284
rect -1544 256 -1516 284
rect -3704 -234 -3676 54
rect -2504 -234 -2476 54
rect -2144 -234 -2116 54
rect -944 -234 -916 54
<< metal4 >>
rect -4320 1014 -4260 1020
rect -4320 726 -4304 1014
rect -4276 726 -4260 1014
rect -4320 720 -4260 726
rect -3360 1014 -3300 1020
rect -3360 726 -3344 1014
rect -3316 726 -3300 1014
rect -3360 720 -3300 726
rect -1320 1014 -1260 1020
rect -1320 726 -1304 1014
rect -1276 726 -1260 1014
rect -1320 720 -1260 726
rect -360 1014 -300 1020
rect -360 726 -344 1014
rect -316 726 -300 1014
rect -360 720 -300 726
rect -4560 524 -4500 540
rect -4560 496 -4544 524
rect -4516 496 -4500 524
rect -4560 480 -4500 496
rect -3960 524 -3900 540
rect -3960 496 -3944 524
rect -3916 496 -3900 524
rect -3960 480 -3900 496
rect -720 524 -660 540
rect -720 496 -704 524
rect -676 496 -660 524
rect -720 480 -660 496
rect -120 524 -60 540
rect -120 496 -104 524
rect -76 496 -60 524
rect -120 480 -60 496
rect -3120 284 -3060 300
rect -3120 256 -3104 284
rect -3076 256 -3060 284
rect -3120 240 -3060 256
rect -2760 284 -2700 300
rect -2760 256 -2744 284
rect -2716 256 -2700 284
rect -2760 240 -2700 256
rect -1920 284 -1860 300
rect -1920 256 -1904 284
rect -1876 256 -1860 284
rect -1920 240 -1860 256
rect -1560 284 -1500 300
rect -1560 256 -1544 284
rect -1516 256 -1500 284
rect -1560 240 -1500 256
rect -3720 54 -3660 60
rect -3720 -234 -3704 54
rect -3676 -234 -3660 54
rect -3720 -240 -3660 -234
rect -2520 54 -2460 60
rect -2520 -234 -2504 54
rect -2476 -234 -2460 54
rect -2520 -240 -2460 -234
rect -2160 54 -2100 60
rect -2160 -234 -2144 54
rect -2116 -234 -2100 54
rect -2160 -240 -2100 -234
rect -960 54 -900 60
rect -960 -234 -944 54
rect -916 -234 -900 54
rect -960 -240 -900 -234
use nauta_cell  nauta_cell_0
timestamp 1665184495
transform 1 0 2460 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_1
timestamp 1665184495
transform 1 0 3060 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_2
timestamp 1665184495
transform 1 0 1860 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_3
timestamp 1665184495
transform 1 0 1260 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_4
timestamp 1665184495
transform 1 0 660 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_5
timestamp 1665184495
transform 1 0 60 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_6
timestamp 1665184495
transform 1 0 -540 0 1 -180
box -3600 -660 -2940 2820
use nauta_cell  nauta_cell_7
timestamp 1665184495
transform 1 0 -1140 0 1 -180
box -3600 -660 -2940 2820
use nauta_edge  nauta_edge_0
timestamp 1665184495
transform -1 0 -3240 0 1 -180
box -3780 -660 -3300 2820
use nauta_edge  nauta_edge_1
timestamp 1665184495
transform 1 0 -1380 0 1 -180
box -3780 -660 -3300 2820
<< labels >>
rlabel metal3 s -5220 240 -5160 300 4 ip
port 1 nsew
rlabel metal3 s -5220 480 -5160 540 4 im
port 2 nsew
rlabel metal3 s -5220 720 -5160 1020 4 op
port 3 nsew
rlabel metal3 s -5220 -240 -5160 60 4 om
port 4 nsew
rlabel metal3 s -5220 2220 -5160 2520 4 vdd
port 5 nsew
rlabel metal3 s -5220 1860 -5160 1920 4 gp
port 6 nsew
rlabel metal3 s -5220 1200 -5160 1260 4 bp
port 7 nsew
rlabel metal3 s -5220 1980 -5160 2040 4 vreg
port 8 nsew
rlabel metal3 s -5220 -840 -5160 -540 4 gnd
port 9 nsew
<< end >>
