magic
tech gf180mcuC
magscale 1 5
timestamp 1665184495
<< metal1 >>
rect -5040 1440 -4980 1500
rect 5160 1440 5220 1500
<< metal2 >>
rect -4440 1254 -4380 1260
rect -4440 966 -4424 1254
rect -4396 966 -4380 1254
rect -4440 960 -4380 966
rect -2040 1254 -1980 1260
rect -2040 966 -2024 1254
rect -1996 966 -1980 1254
rect -2040 960 -1980 966
rect -240 1254 -180 1260
rect -240 966 -224 1254
rect -196 966 -180 1254
rect -240 960 -180 966
rect 360 1254 420 1260
rect 360 966 376 1254
rect 404 966 420 1254
rect 360 960 420 966
rect 2160 1254 2220 1260
rect 2160 966 2176 1254
rect 2204 966 2220 1254
rect 2160 960 2220 966
rect 4560 1254 4620 1260
rect 4560 966 4576 1254
rect 4604 966 4620 1254
rect 4560 960 4620 966
rect -3240 524 -3180 540
rect -3240 496 -3224 524
rect -3196 496 -3180 524
rect -3240 480 -3180 496
rect -2640 524 -2580 540
rect -2640 496 -2624 524
rect -2596 496 -2580 524
rect -2640 480 -2580 496
rect 2760 524 2820 540
rect 2760 496 2776 524
rect 2804 496 2820 524
rect 2760 480 2820 496
rect 3360 524 3420 540
rect 3360 496 3376 524
rect 3404 496 3420 524
rect 3360 480 3420 496
rect -3840 54 -3780 60
rect -3840 -234 -3824 54
rect -3796 -234 -3780 54
rect -3840 -240 -3780 -234
rect -1440 54 -1380 60
rect -1440 -234 -1424 54
rect -1396 -234 -1380 54
rect -1440 -240 -1380 -234
rect -840 54 -780 60
rect -840 -234 -824 54
rect -796 -234 -780 54
rect -840 -240 -780 -234
rect 960 54 1020 60
rect 960 -234 976 54
rect 1004 -234 1020 54
rect 960 -240 1020 -234
rect 1560 54 1620 60
rect 1560 -234 1576 54
rect 1604 -234 1620 54
rect 1560 -240 1620 -234
rect 3960 54 4020 60
rect 3960 -234 3976 54
rect 4004 -234 4020 54
rect 3960 -240 4020 -234
<< via2 >>
rect -4424 966 -4396 1254
rect -2024 966 -1996 1254
rect -224 966 -196 1254
rect 376 966 404 1254
rect 2176 966 2204 1254
rect 4576 966 4604 1254
rect -3224 496 -3196 524
rect -2624 496 -2596 524
rect 2776 496 2804 524
rect 3376 496 3404 524
rect -3824 -234 -3796 54
rect -1424 -234 -1396 54
rect -824 -234 -796 54
rect 976 -234 1004 54
rect 1576 -234 1604 54
rect 3976 -234 4004 54
<< metal3 >>
rect -5220 2460 -5160 2760
rect -5220 2190 -5160 2280
rect -5220 2100 -5160 2160
rect -5220 1440 -2280 1500
rect 2460 1440 5340 1500
rect -5220 960 -5160 1260
rect -4440 1254 -4380 1260
rect -4440 966 -4424 1254
rect -4396 966 -4380 1254
rect -4440 960 -4380 966
rect -2160 1254 -2100 1260
rect -2160 966 -2144 1254
rect -2116 966 -2100 1254
rect -2160 960 -2100 966
rect -2040 1254 -1980 1260
rect -2040 966 -2024 1254
rect -1996 966 -1980 1254
rect -2040 960 -1980 966
rect -1320 1254 -1260 1260
rect -1320 966 -1304 1254
rect -1276 966 -1260 1254
rect -1320 960 -1260 966
rect -240 1254 -180 1260
rect -240 966 -224 1254
rect -196 966 -180 1254
rect -240 960 -180 966
rect 360 1254 420 1260
rect 360 966 376 1254
rect 404 966 420 1254
rect 360 960 420 966
rect 1440 1254 1500 1260
rect 1440 966 1456 1254
rect 1484 966 1500 1254
rect 1440 960 1500 966
rect 2160 1254 2220 1260
rect 2160 966 2176 1254
rect 2204 966 2220 1254
rect 2160 960 2220 966
rect 2280 1254 2340 1260
rect 2280 966 2296 1254
rect 2324 966 2340 1254
rect 2280 960 2340 966
rect 4560 1254 4620 1260
rect 4560 966 4576 1254
rect 4604 966 4620 1254
rect 4560 960 4620 966
rect -5220 720 -5160 780
rect -4560 764 -4500 780
rect -4560 736 -4544 764
rect -4516 736 -4500 764
rect -4560 720 -4500 736
rect -2520 764 -2460 780
rect -2520 736 -2504 764
rect -2476 736 -2460 764
rect -2520 720 -2460 736
rect -120 764 -60 780
rect -120 736 -104 764
rect -76 736 -60 764
rect -120 720 -60 736
rect 240 764 300 780
rect 240 736 256 764
rect 284 736 300 764
rect 240 720 300 736
rect 2640 764 2700 780
rect 2640 736 2656 764
rect 2684 736 2700 764
rect 2640 720 2700 736
rect 4680 764 4740 780
rect 4680 736 4696 764
rect 4724 736 4740 764
rect 4680 720 4740 736
rect -5220 480 -5160 540
rect -4320 524 -4260 540
rect -4320 496 -4304 524
rect -4276 496 -4260 524
rect -4320 480 -4260 496
rect -3960 524 -3900 540
rect -3960 496 -3944 524
rect -3916 496 -3900 524
rect -3960 480 -3900 496
rect -3240 524 -3180 540
rect -3240 496 -3224 524
rect -3196 496 -3180 524
rect -3240 480 -3180 496
rect -3120 524 -3060 540
rect -3120 496 -3104 524
rect -3076 496 -3060 524
rect -3120 480 -3060 496
rect -2760 524 -2700 540
rect -2760 496 -2744 524
rect -2716 496 -2700 524
rect -2760 480 -2700 496
rect -2640 524 -2580 540
rect -2640 496 -2624 524
rect -2596 496 -2580 524
rect -2640 480 -2580 496
rect -720 524 -660 540
rect -720 496 -704 524
rect -676 496 -660 524
rect -720 480 -660 496
rect -360 524 -300 540
rect -360 496 -344 524
rect -316 496 -300 524
rect -360 480 -300 496
rect 480 524 540 540
rect 480 496 496 524
rect 524 496 540 524
rect 480 480 540 496
rect 840 524 900 540
rect 840 496 856 524
rect 884 496 900 524
rect 840 480 900 496
rect 2760 524 2820 540
rect 2760 496 2776 524
rect 2804 496 2820 524
rect 2760 480 2820 496
rect 2880 524 2940 540
rect 2880 496 2896 524
rect 2924 496 2940 524
rect 2880 480 2940 496
rect 3240 524 3300 540
rect 3240 496 3256 524
rect 3284 496 3300 524
rect 3240 480 3300 496
rect 3360 524 3420 540
rect 3360 496 3376 524
rect 3404 496 3420 524
rect 3360 480 3420 496
rect 4080 524 4140 540
rect 4080 496 4096 524
rect 4124 496 4140 524
rect 4080 480 4140 496
rect 4440 524 4500 540
rect 4440 496 4456 524
rect 4484 496 4500 524
rect 4440 480 4500 496
rect -5220 240 -5160 300
rect -3720 284 -3660 300
rect -3720 256 -3704 284
rect -3676 256 -3660 284
rect -3720 240 -3660 256
rect -3360 284 -3300 300
rect -3360 256 -3344 284
rect -3316 256 -3300 284
rect -3360 240 -3300 256
rect -960 284 -900 300
rect -960 256 -944 284
rect -916 256 -900 284
rect -960 240 -900 256
rect 1080 284 1140 300
rect 1080 256 1096 284
rect 1124 256 1140 284
rect 1080 240 1140 256
rect 3480 284 3540 300
rect 3480 256 3496 284
rect 3524 256 3540 284
rect 3480 240 3540 256
rect 3840 284 3900 300
rect 3840 256 3856 284
rect 3884 256 3900 284
rect 3840 240 3900 256
rect -5220 -240 -5160 60
rect -3840 54 -3780 60
rect -3840 -234 -3824 54
rect -3796 -234 -3780 54
rect -3840 -240 -3780 -234
rect -1920 54 -1860 60
rect -1920 -234 -1904 54
rect -1876 -234 -1860 54
rect -1920 -240 -1860 -234
rect -1560 54 -1500 60
rect -1560 -234 -1544 54
rect -1516 -234 -1500 54
rect -1560 -240 -1500 -234
rect -1440 54 -1380 60
rect -1440 -234 -1424 54
rect -1396 -234 -1380 54
rect -1440 -240 -1380 -234
rect -840 54 -780 60
rect -840 -234 -824 54
rect -796 -234 -780 54
rect -840 -240 -780 -234
rect 960 54 1020 60
rect 960 -234 976 54
rect 1004 -234 1020 54
rect 960 -240 1020 -234
rect 1560 54 1620 60
rect 1560 -234 1576 54
rect 1604 -234 1620 54
rect 1560 -240 1620 -234
rect 1680 54 1740 60
rect 1680 -234 1696 54
rect 1724 -234 1740 54
rect 1680 -240 1740 -234
rect 2040 54 2100 60
rect 2040 -234 2056 54
rect 2084 -234 2100 54
rect 2040 -240 2100 -234
rect 3960 54 4020 60
rect 3960 -234 3976 54
rect 4004 -234 4020 54
rect 3960 -240 4020 -234
rect -5220 -840 -5160 -540
<< via3 >>
rect -2144 966 -2116 1254
rect -1304 966 -1276 1254
rect 1456 966 1484 1254
rect 2296 966 2324 1254
rect -4544 736 -4516 764
rect -2504 736 -2476 764
rect -104 736 -76 764
rect 256 736 284 764
rect 2656 736 2684 764
rect 4696 736 4724 764
rect -4304 496 -4276 524
rect -3944 496 -3916 524
rect -3104 496 -3076 524
rect -2744 496 -2716 524
rect -704 496 -676 524
rect -344 496 -316 524
rect 496 496 524 524
rect 856 496 884 524
rect 2896 496 2924 524
rect 3256 496 3284 524
rect 4096 496 4124 524
rect 4456 496 4484 524
rect -3704 256 -3676 284
rect -3344 256 -3316 284
rect -944 256 -916 284
rect 1096 256 1124 284
rect 3496 256 3524 284
rect 3856 256 3884 284
rect -1904 -234 -1876 54
rect -1544 -234 -1516 54
rect 1696 -234 1724 54
rect 2056 -234 2084 54
<< metal4 >>
rect -2160 1254 -2100 1260
rect -2160 966 -2144 1254
rect -2116 966 -2100 1254
rect -2160 960 -2100 966
rect -1320 1254 -1260 1260
rect -1320 966 -1304 1254
rect -1276 966 -1260 1254
rect -1320 960 -1260 966
rect 1440 1254 1500 1260
rect 1440 966 1456 1254
rect 1484 966 1500 1254
rect 1440 960 1500 966
rect 2280 1254 2340 1260
rect 2280 966 2296 1254
rect 2324 966 2340 1254
rect 2280 960 2340 966
rect -4560 764 -4500 780
rect -4560 736 -4544 764
rect -4516 736 -4500 764
rect -4560 720 -4500 736
rect -2520 764 -2460 780
rect -2520 736 -2504 764
rect -2476 736 -2460 764
rect -2520 720 -2460 736
rect -120 764 -60 780
rect -120 736 -104 764
rect -76 736 -60 764
rect -120 720 -60 736
rect 240 764 300 780
rect 240 736 256 764
rect 284 736 300 764
rect 240 720 300 736
rect 2640 764 2700 780
rect 2640 736 2656 764
rect 2684 736 2700 764
rect 2640 720 2700 736
rect 4680 764 4740 780
rect 4680 736 4696 764
rect 4724 736 4740 764
rect 4680 720 4740 736
rect -4320 524 -4260 540
rect -4320 496 -4304 524
rect -4276 496 -4260 524
rect -4320 480 -4260 496
rect -3960 524 -3900 540
rect -3960 496 -3944 524
rect -3916 496 -3900 524
rect -3960 480 -3900 496
rect -3120 524 -3060 540
rect -3120 496 -3104 524
rect -3076 496 -3060 524
rect -3120 480 -3060 496
rect -2760 524 -2700 540
rect -2760 496 -2744 524
rect -2716 496 -2700 524
rect -2760 480 -2700 496
rect -720 524 -660 540
rect -720 496 -704 524
rect -676 496 -660 524
rect -720 480 -660 496
rect -360 524 -300 540
rect -360 496 -344 524
rect -316 496 -300 524
rect -360 480 -300 496
rect 480 524 540 540
rect 480 496 496 524
rect 524 496 540 524
rect 480 480 540 496
rect 840 524 900 540
rect 840 496 856 524
rect 884 496 900 524
rect 840 480 900 496
rect 2880 524 2940 540
rect 2880 496 2896 524
rect 2924 496 2940 524
rect 2880 480 2940 496
rect 3240 524 3300 540
rect 3240 496 3256 524
rect 3284 496 3300 524
rect 3240 480 3300 496
rect 4080 524 4140 540
rect 4080 496 4096 524
rect 4124 496 4140 524
rect 4080 480 4140 496
rect 4440 524 4500 540
rect 4440 496 4456 524
rect 4484 496 4500 524
rect 4440 480 4500 496
rect -3720 284 -3660 300
rect -3720 256 -3704 284
rect -3676 256 -3660 284
rect -3720 240 -3660 256
rect -3360 284 -3300 300
rect -3360 256 -3344 284
rect -3316 256 -3300 284
rect -3360 240 -3300 256
rect -960 284 -900 300
rect -960 256 -944 284
rect -916 256 -900 284
rect -960 240 -900 256
rect 1080 284 1140 300
rect 1080 256 1096 284
rect 1124 256 1140 284
rect 1080 240 1140 256
rect 3480 284 3540 300
rect 3480 256 3496 284
rect 3524 256 3540 284
rect 3480 240 3540 256
rect 3840 284 3900 300
rect 3840 256 3856 284
rect 3884 256 3900 284
rect 3840 240 3900 256
rect -1920 54 -1860 60
rect -1920 -234 -1904 54
rect -1876 -234 -1860 54
rect -1920 -240 -1860 -234
rect -1560 54 -1500 60
rect -1560 -234 -1544 54
rect -1516 -234 -1500 54
rect -1560 -240 -1500 -234
rect 1680 54 1740 60
rect 1680 -234 1696 54
rect 1724 -234 1740 54
rect 1680 -240 1740 -234
rect 2040 54 2100 60
rect 2040 -234 2056 54
rect 2084 -234 2100 54
rect 2040 -240 2100 -234
use barthnauta_cell  barthnauta_cell_0
timestamp 1665184495
transform -1 0 1320 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_1
timestamp 1665184495
transform -1 0 720 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_2
timestamp 1665184495
transform -1 0 120 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_3
timestamp 1665184495
transform -1 0 -480 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_4
timestamp 1665184495
transform -1 0 -1080 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_5
timestamp 1665184495
transform -1 0 -1680 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_6
timestamp 1665184495
transform -1 0 -2280 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_7
timestamp 1665184495
transform -1 0 -2880 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_8
timestamp 1665184495
transform 1 0 3060 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_9
timestamp 1665184495
transform 1 0 2460 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_10
timestamp 1665184495
transform 1 0 1860 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_11
timestamp 1665184495
transform 1 0 1260 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_12
timestamp 1665184495
transform 1 0 660 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_13
timestamp 1665184495
transform 1 0 60 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_14
timestamp 1665184495
transform 1 0 -540 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_cell  barthnauta_cell_15
timestamp 1665184495
transform 1 0 -1140 0 1 -180
box -3600 -660 -2940 3060
use barthnauta_edge  barthnauta_edge_0
timestamp 1665184495
transform -1 0 1560 0 1 -180
box -3780 -660 -3300 3060
use barthnauta_edge  barthnauta_edge_1
timestamp 1665184495
transform 1 0 -1380 0 1 -180
box -3780 -660 -3300 3060
<< labels >>
rlabel metal3 s -5190 510 -5190 510 4 x
rlabel metal3 s -5220 240 -5160 300 4 ip
port 1 nsew
rlabel metal3 s -5220 720 -5160 780 4 im
port 2 nsew
rlabel metal3 s -5220 960 -5160 1260 4 op
port 3 nsew
rlabel metal3 s -5220 -240 -5160 60 4 om
port 4 nsew
rlabel metal3 s -5220 2460 -5160 2760 4 vdd
port 5 nsew
rlabel metal3 s -5220 2100 -5160 2160 4 gp
port 6 nsew
rlabel metal3 s -5220 1440 -5160 1500 4 bp
port 7 nsew
rlabel metal3 s -5220 2220 -5160 2280 4 vreg
port 8 nsew
rlabel metal3 s -5220 -840 -5160 -540 4 gnd
port 9 nsew
<< end >>
