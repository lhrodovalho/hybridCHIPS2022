magic
tech gf180mcuC
timestamp 1663271470
<< nwell >>
rect -720 474 -588 594
rect -720 318 -588 450
<< nmos >>
rect -696 -108 -684 -72
rect -672 -108 -660 -72
rect -648 -108 -636 -72
rect -624 -108 -612 -72
<< pmos >>
rect -696 372 -684 402
rect -672 372 -660 402
rect -648 372 -636 402
rect -624 372 -612 402
<< mvpmos >>
rect -696 528 -684 564
rect -672 528 -660 564
rect -648 528 -636 564
rect -624 528 -612 564
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
<< pdiff >>
rect -708 393 -696 402
rect -708 387 -705 393
rect -699 387 -696 393
rect -708 381 -696 387
rect -708 375 -705 381
rect -699 375 -696 381
rect -708 372 -696 375
rect -684 393 -672 402
rect -684 387 -681 393
rect -675 387 -672 393
rect -684 381 -672 387
rect -684 375 -681 381
rect -675 375 -672 381
rect -684 372 -672 375
rect -660 393 -648 402
rect -660 387 -657 393
rect -651 387 -648 393
rect -660 381 -648 387
rect -660 375 -657 381
rect -651 375 -648 381
rect -660 372 -648 375
rect -636 393 -624 402
rect -636 387 -633 393
rect -627 387 -624 393
rect -636 381 -624 387
rect -636 375 -633 381
rect -627 375 -624 381
rect -636 372 -624 375
rect -612 393 -600 402
rect -612 387 -609 393
rect -603 387 -600 393
rect -612 381 -600 387
rect -612 375 -609 381
rect -603 375 -600 381
rect -612 372 -600 375
<< mvpdiff >>
rect -708 561 -696 564
rect -708 555 -705 561
rect -699 555 -696 561
rect -708 549 -696 555
rect -708 543 -705 549
rect -699 543 -696 549
rect -708 537 -696 543
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 528 -696 531
rect -684 561 -672 564
rect -684 555 -681 561
rect -675 555 -672 561
rect -684 549 -672 555
rect -684 543 -681 549
rect -675 543 -672 549
rect -684 537 -672 543
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 528 -672 531
rect -660 561 -648 564
rect -660 555 -657 561
rect -651 555 -648 561
rect -660 549 -648 555
rect -660 543 -657 549
rect -651 543 -648 549
rect -660 537 -648 543
rect -660 531 -657 537
rect -651 531 -648 537
rect -660 528 -648 531
rect -636 561 -624 564
rect -636 555 -633 561
rect -627 555 -624 561
rect -636 549 -624 555
rect -636 543 -633 549
rect -627 543 -624 549
rect -636 537 -624 543
rect -636 531 -633 537
rect -627 531 -624 537
rect -636 528 -624 531
rect -612 561 -600 564
rect -612 555 -609 561
rect -603 555 -600 561
rect -612 549 -600 555
rect -612 543 -609 549
rect -603 543 -600 549
rect -612 537 -600 543
rect -612 531 -609 537
rect -603 531 -600 537
rect -612 528 -600 531
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -633 -81 -627 -75
rect -633 -93 -627 -87
rect -633 -105 -627 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
<< pdiffc >>
rect -705 387 -699 393
rect -705 375 -699 381
rect -681 387 -675 393
rect -681 375 -675 381
rect -657 387 -651 393
rect -657 375 -651 381
rect -633 387 -627 393
rect -633 375 -627 381
rect -609 387 -603 393
rect -609 375 -603 381
<< mvpdiffc >>
rect -705 555 -699 561
rect -705 543 -699 549
rect -705 531 -699 537
rect -681 555 -675 561
rect -681 543 -675 549
rect -681 531 -675 537
rect -657 555 -651 561
rect -657 543 -651 549
rect -657 531 -651 537
rect -633 555 -627 561
rect -633 543 -627 549
rect -633 531 -627 537
rect -609 555 -603 561
rect -609 543 -603 549
rect -609 531 -603 537
<< psubdiff >>
rect -720 609 -588 612
rect -720 603 -717 609
rect -711 603 -705 609
rect -699 603 -693 609
rect -687 603 -681 609
rect -675 603 -669 609
rect -663 603 -657 609
rect -651 603 -645 609
rect -639 603 -633 609
rect -627 603 -621 609
rect -615 603 -609 609
rect -603 603 -597 609
rect -591 603 -588 609
rect -720 600 -588 603
rect -720 465 -588 468
rect -720 459 -717 465
rect -711 459 -705 465
rect -699 459 -693 465
rect -687 459 -681 465
rect -675 459 -669 465
rect -663 459 -657 465
rect -651 459 -645 465
rect -639 459 -633 465
rect -627 459 -621 465
rect -615 459 -609 465
rect -603 459 -597 465
rect -591 459 -588 465
rect -720 456 -588 459
rect -720 309 -588 312
rect -720 303 -717 309
rect -711 303 -705 309
rect -699 303 -693 309
rect -687 303 -681 309
rect -675 303 -669 309
rect -663 303 -657 309
rect -651 303 -645 309
rect -639 303 -633 309
rect -627 303 -621 309
rect -615 303 -609 309
rect -603 303 -597 309
rect -591 303 -588 309
rect -720 300 -588 303
rect -720 213 -588 216
rect -720 207 -717 213
rect -711 207 -705 213
rect -699 207 -693 213
rect -687 207 -681 213
rect -675 207 -669 213
rect -663 207 -657 213
rect -651 207 -645 213
rect -639 207 -633 213
rect -627 207 -621 213
rect -615 207 -609 213
rect -603 207 -597 213
rect -591 207 -588 213
rect -720 204 -588 207
rect -720 165 -588 168
rect -720 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -657 165
rect -651 159 -645 165
rect -639 159 -633 165
rect -627 159 -621 165
rect -615 159 -609 165
rect -603 159 -597 165
rect -591 159 -588 165
rect -720 156 -588 159
rect -720 117 -588 120
rect -720 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -657 117
rect -651 111 -645 117
rect -639 111 -633 117
rect -627 111 -621 117
rect -615 111 -609 117
rect -603 111 -597 117
rect -591 111 -588 117
rect -720 108 -588 111
rect -720 69 -588 72
rect -720 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -657 69
rect -651 63 -645 69
rect -639 63 -633 69
rect -627 63 -621 69
rect -615 63 -609 69
rect -603 63 -597 69
rect -591 63 -588 69
rect -720 60 -588 63
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< nsubdiff >>
rect -708 441 -600 444
rect -708 435 -705 441
rect -699 435 -693 441
rect -687 435 -681 441
rect -675 435 -669 441
rect -663 435 -657 441
rect -651 435 -645 441
rect -639 435 -633 441
rect -627 435 -621 441
rect -615 435 -609 441
rect -603 435 -600 441
rect -708 432 -600 435
rect -708 333 -600 336
rect -708 327 -705 333
rect -699 327 -693 333
rect -687 327 -681 333
rect -675 327 -669 333
rect -663 327 -657 333
rect -651 327 -645 333
rect -639 327 -633 333
rect -627 327 -621 333
rect -615 327 -609 333
rect -603 327 -600 333
rect -708 324 -600 327
<< mvnsubdiff >>
rect -708 585 -600 588
rect -708 579 -705 585
rect -699 579 -693 585
rect -687 579 -681 585
rect -675 579 -669 585
rect -663 579 -657 585
rect -651 579 -645 585
rect -639 579 -633 585
rect -627 579 -621 585
rect -615 579 -609 585
rect -603 579 -600 585
rect -708 576 -600 579
rect -708 489 -600 492
rect -708 483 -705 489
rect -699 483 -693 489
rect -687 483 -681 489
rect -675 483 -669 489
rect -663 483 -657 489
rect -651 483 -645 489
rect -639 483 -633 489
rect -627 483 -621 489
rect -615 483 -609 489
rect -603 483 -600 489
rect -708 480 -600 483
<< psubdiffcont >>
rect -717 603 -711 609
rect -705 603 -699 609
rect -693 603 -687 609
rect -681 603 -675 609
rect -669 603 -663 609
rect -657 603 -651 609
rect -645 603 -639 609
rect -633 603 -627 609
rect -621 603 -615 609
rect -609 603 -603 609
rect -597 603 -591 609
rect -717 459 -711 465
rect -705 459 -699 465
rect -693 459 -687 465
rect -681 459 -675 465
rect -669 459 -663 465
rect -657 459 -651 465
rect -645 459 -639 465
rect -633 459 -627 465
rect -621 459 -615 465
rect -609 459 -603 465
rect -597 459 -591 465
rect -717 303 -711 309
rect -705 303 -699 309
rect -693 303 -687 309
rect -681 303 -675 309
rect -669 303 -663 309
rect -657 303 -651 309
rect -645 303 -639 309
rect -633 303 -627 309
rect -621 303 -615 309
rect -609 303 -603 309
rect -597 303 -591 309
rect -717 207 -711 213
rect -705 207 -699 213
rect -693 207 -687 213
rect -681 207 -675 213
rect -669 207 -663 213
rect -657 207 -651 213
rect -645 207 -639 213
rect -633 207 -627 213
rect -621 207 -615 213
rect -609 207 -603 213
rect -597 207 -591 213
rect -717 159 -711 165
rect -705 159 -699 165
rect -693 159 -687 165
rect -681 159 -675 165
rect -669 159 -663 165
rect -657 159 -651 165
rect -645 159 -639 165
rect -633 159 -627 165
rect -621 159 -615 165
rect -609 159 -603 165
rect -597 159 -591 165
rect -717 111 -711 117
rect -705 111 -699 117
rect -693 111 -687 117
rect -681 111 -675 117
rect -669 111 -663 117
rect -657 111 -651 117
rect -645 111 -639 117
rect -633 111 -627 117
rect -621 111 -615 117
rect -609 111 -603 117
rect -597 111 -591 117
rect -717 63 -711 69
rect -705 63 -699 69
rect -693 63 -687 69
rect -681 63 -675 69
rect -669 63 -663 69
rect -657 63 -651 69
rect -645 63 -639 69
rect -633 63 -627 69
rect -621 63 -615 69
rect -609 63 -603 69
rect -597 63 -591 69
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -657 -33 -651 -27
rect -645 -33 -639 -27
rect -633 -33 -627 -27
rect -621 -33 -615 -27
rect -609 -33 -603 -27
rect -597 -33 -591 -27
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
rect -657 -129 -651 -123
rect -645 -129 -639 -123
rect -633 -129 -627 -123
rect -621 -129 -615 -123
rect -609 -129 -603 -123
rect -597 -129 -591 -123
<< nsubdiffcont >>
rect -705 435 -699 441
rect -693 435 -687 441
rect -681 435 -675 441
rect -669 435 -663 441
rect -657 435 -651 441
rect -645 435 -639 441
rect -633 435 -627 441
rect -621 435 -615 441
rect -609 435 -603 441
rect -705 327 -699 333
rect -693 327 -687 333
rect -681 327 -675 333
rect -669 327 -663 333
rect -657 327 -651 333
rect -645 327 -639 333
rect -633 327 -627 333
rect -621 327 -615 333
rect -609 327 -603 333
<< mvnsubdiffcont >>
rect -705 579 -699 585
rect -693 579 -687 585
rect -681 579 -675 585
rect -669 579 -663 585
rect -657 579 -651 585
rect -645 579 -639 585
rect -633 579 -627 585
rect -621 579 -615 585
rect -609 579 -603 585
rect -705 483 -699 489
rect -693 483 -687 489
rect -681 483 -675 489
rect -669 483 -663 489
rect -657 483 -651 489
rect -645 483 -639 489
rect -633 483 -627 489
rect -621 483 -615 489
rect -609 483 -603 489
<< polysilicon >>
rect -696 564 -684 570
rect -672 564 -660 570
rect -648 564 -636 570
rect -624 564 -612 570
rect -696 516 -684 528
rect -672 516 -660 528
rect -648 516 -636 528
rect -624 516 -612 528
rect -696 513 -612 516
rect -696 507 -693 513
rect -687 507 -681 513
rect -675 507 -669 513
rect -663 507 -657 513
rect -651 507 -645 513
rect -639 507 -633 513
rect -627 507 -621 513
rect -615 507 -612 513
rect -696 504 -612 507
rect -696 402 -684 408
rect -672 402 -660 408
rect -648 402 -636 408
rect -624 402 -612 408
rect -696 360 -684 372
rect -672 360 -660 372
rect -696 357 -660 360
rect -696 351 -693 357
rect -687 351 -681 357
rect -675 351 -669 357
rect -663 351 -660 357
rect -696 348 -660 351
rect -648 360 -636 372
rect -624 360 -612 372
rect -648 357 -612 360
rect -648 351 -645 357
rect -639 351 -633 357
rect -627 351 -621 357
rect -615 351 -612 357
rect -648 348 -612 351
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -696 -72 -684 -60
rect -672 -72 -660 -60
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -648 -72 -636 -60
rect -624 -72 -612 -60
rect -696 -114 -684 -108
rect -672 -114 -660 -108
rect -648 -114 -636 -108
rect -624 -114 -612 -108
<< polycontact >>
rect -693 507 -687 513
rect -681 507 -675 513
rect -669 507 -663 513
rect -657 507 -651 513
rect -645 507 -639 513
rect -633 507 -627 513
rect -621 507 -615 513
rect -693 351 -687 357
rect -681 351 -675 357
rect -669 351 -663 357
rect -645 351 -639 357
rect -633 351 -627 357
rect -621 351 -615 357
rect -693 -57 -687 -51
rect -681 -57 -675 -51
rect -669 -57 -663 -51
rect -645 -57 -639 -51
rect -633 -57 -627 -51
rect -621 -57 -615 -51
<< metal1 >>
rect -720 609 -588 612
rect -720 603 -717 609
rect -711 603 -705 609
rect -699 603 -693 609
rect -687 603 -681 609
rect -675 603 -669 609
rect -663 603 -657 609
rect -651 603 -645 609
rect -639 603 -633 609
rect -627 603 -621 609
rect -615 603 -609 609
rect -603 603 -597 609
rect -591 603 -588 609
rect -720 600 -588 603
rect -720 585 -588 588
rect -720 579 -705 585
rect -699 579 -693 585
rect -687 579 -681 585
rect -675 579 -669 585
rect -663 579 -657 585
rect -651 579 -645 585
rect -639 579 -633 585
rect -627 579 -621 585
rect -615 579 -609 585
rect -603 579 -588 585
rect -720 576 -588 579
rect -708 561 -696 564
rect -708 555 -705 561
rect -699 555 -696 561
rect -708 549 -696 555
rect -708 543 -705 549
rect -699 543 -696 549
rect -708 537 -696 543
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 528 -696 531
rect -684 561 -672 564
rect -684 555 -681 561
rect -675 555 -672 561
rect -684 549 -672 555
rect -684 543 -681 549
rect -675 543 -672 549
rect -684 537 -672 543
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 528 -672 531
rect -660 561 -648 564
rect -660 555 -657 561
rect -651 555 -648 561
rect -660 549 -648 555
rect -660 543 -657 549
rect -651 543 -648 549
rect -660 537 -648 543
rect -660 531 -657 537
rect -651 531 -648 537
rect -660 528 -648 531
rect -636 561 -624 564
rect -636 555 -633 561
rect -627 555 -624 561
rect -636 549 -624 555
rect -636 543 -633 549
rect -627 543 -624 549
rect -636 537 -624 543
rect -636 531 -633 537
rect -627 531 -624 537
rect -636 528 -624 531
rect -612 561 -600 564
rect -612 555 -609 561
rect -603 555 -600 561
rect -612 549 -600 555
rect -612 543 -609 549
rect -603 543 -600 549
rect -612 537 -600 543
rect -612 531 -609 537
rect -603 531 -600 537
rect -612 528 -600 531
rect -696 513 -612 516
rect -696 507 -693 513
rect -687 507 -681 513
rect -675 507 -669 513
rect -663 507 -657 513
rect -651 507 -645 513
rect -639 507 -633 513
rect -627 507 -621 513
rect -615 507 -612 513
rect -696 504 -612 507
rect -720 489 -588 492
rect -720 483 -705 489
rect -699 483 -693 489
rect -687 483 -681 489
rect -675 483 -669 489
rect -663 483 -657 489
rect -651 483 -645 489
rect -639 483 -633 489
rect -627 483 -621 489
rect -615 483 -609 489
rect -603 483 -588 489
rect -720 480 -588 483
rect -720 465 -588 468
rect -720 459 -717 465
rect -711 459 -705 465
rect -699 459 -693 465
rect -687 459 -681 465
rect -675 459 -669 465
rect -663 459 -657 465
rect -651 459 -645 465
rect -639 459 -633 465
rect -627 459 -621 465
rect -615 459 -609 465
rect -603 459 -597 465
rect -591 459 -588 465
rect -720 456 -588 459
rect -720 441 -588 444
rect -720 435 -705 441
rect -699 435 -693 441
rect -687 435 -681 441
rect -675 435 -669 441
rect -663 435 -657 441
rect -651 435 -645 441
rect -639 435 -633 441
rect -627 435 -621 441
rect -615 435 -609 441
rect -603 435 -588 441
rect -720 432 -588 435
rect -708 417 -600 420
rect -708 411 -705 417
rect -699 411 -657 417
rect -651 411 -609 417
rect -603 411 -600 417
rect -708 408 -600 411
rect -708 405 -696 408
rect -708 399 -705 405
rect -699 399 -696 405
rect -660 405 -648 408
rect -708 393 -696 399
rect -708 387 -705 393
rect -699 387 -696 393
rect -708 381 -696 387
rect -708 375 -705 381
rect -699 375 -696 381
rect -708 372 -696 375
rect -684 393 -672 402
rect -684 387 -681 393
rect -675 387 -672 393
rect -684 381 -672 387
rect -684 375 -681 381
rect -675 375 -672 381
rect -684 372 -672 375
rect -660 399 -657 405
rect -651 399 -648 405
rect -612 405 -600 408
rect -660 393 -648 399
rect -660 387 -657 393
rect -651 387 -648 393
rect -660 381 -648 387
rect -660 375 -657 381
rect -651 375 -648 381
rect -660 372 -648 375
rect -636 393 -624 402
rect -636 387 -633 393
rect -627 387 -624 393
rect -636 381 -624 387
rect -636 375 -633 381
rect -627 375 -624 381
rect -636 372 -624 375
rect -612 399 -609 405
rect -603 399 -600 405
rect -612 393 -600 399
rect -612 387 -609 393
rect -603 387 -600 393
rect -612 381 -600 387
rect -612 375 -609 381
rect -603 375 -600 381
rect -612 372 -600 375
rect -696 357 -660 360
rect -696 351 -693 357
rect -687 351 -681 357
rect -675 351 -669 357
rect -663 351 -660 357
rect -696 348 -660 351
rect -648 357 -612 360
rect -648 351 -645 357
rect -639 351 -633 357
rect -627 351 -621 357
rect -615 351 -612 357
rect -648 348 -612 351
rect -720 333 -588 336
rect -720 327 -705 333
rect -699 327 -693 333
rect -687 327 -681 333
rect -675 327 -669 333
rect -663 327 -657 333
rect -651 327 -645 333
rect -639 327 -633 333
rect -627 327 -621 333
rect -615 327 -609 333
rect -603 327 -588 333
rect -720 324 -588 327
rect -720 309 -588 312
rect -720 303 -717 309
rect -711 303 -705 309
rect -699 303 -693 309
rect -687 303 -681 309
rect -675 303 -669 309
rect -663 303 -657 309
rect -651 303 -645 309
rect -639 303 -633 309
rect -627 303 -621 309
rect -615 303 -609 309
rect -603 303 -597 309
rect -591 303 -588 309
rect -720 300 -588 303
rect -720 213 -588 216
rect -720 207 -717 213
rect -711 207 -705 213
rect -699 207 -693 213
rect -687 207 -681 213
rect -675 207 -669 213
rect -663 207 -657 213
rect -651 207 -645 213
rect -639 207 -633 213
rect -627 207 -621 213
rect -615 207 -609 213
rect -603 207 -597 213
rect -591 207 -588 213
rect -720 204 -588 207
rect -720 165 -588 168
rect -720 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -657 165
rect -651 159 -645 165
rect -639 159 -633 165
rect -627 159 -621 165
rect -615 159 -609 165
rect -603 159 -597 165
rect -591 159 -588 165
rect -720 156 -588 159
rect -720 117 -588 120
rect -720 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -657 117
rect -651 111 -645 117
rect -639 111 -633 117
rect -627 111 -621 117
rect -615 111 -609 117
rect -603 111 -597 117
rect -591 111 -588 117
rect -720 108 -588 111
rect -720 69 -588 72
rect -720 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -657 69
rect -651 63 -645 69
rect -639 63 -633 69
rect -627 63 -621 69
rect -615 63 -609 69
rect -603 63 -597 69
rect -591 63 -588 69
rect -720 60 -588 63
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< via1 >>
rect -705 579 -699 585
rect -657 579 -651 585
rect -609 579 -603 585
rect -705 555 -699 561
rect -705 543 -699 549
rect -705 531 -699 537
rect -681 555 -675 561
rect -681 543 -675 549
rect -681 531 -675 537
rect -657 555 -651 561
rect -657 543 -651 549
rect -657 531 -651 537
rect -633 555 -627 561
rect -633 543 -627 549
rect -633 531 -627 537
rect -609 555 -603 561
rect -609 543 -603 549
rect -609 531 -603 537
rect -657 507 -651 513
rect -705 411 -699 417
rect -657 411 -651 417
rect -609 411 -603 417
rect -705 399 -699 405
rect -705 387 -699 393
rect -705 375 -699 381
rect -681 387 -675 393
rect -681 375 -675 381
rect -657 399 -651 405
rect -633 387 -627 393
rect -633 375 -627 381
rect -609 399 -603 405
rect -609 387 -603 393
rect -609 375 -603 381
rect -681 351 -675 357
rect -633 351 -627 357
rect -705 327 -699 333
rect -609 327 -603 333
rect -705 303 -699 309
rect -609 303 -603 309
rect -705 207 -699 213
rect -609 207 -603 213
rect -705 159 -699 165
rect -609 159 -603 165
rect -705 111 -699 117
rect -609 111 -603 117
rect -705 63 -699 69
rect -609 63 -603 69
rect -705 -33 -699 -27
rect -609 -33 -603 -27
rect -681 -57 -675 -51
rect -633 -57 -627 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal2 >>
rect -708 585 -696 588
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 561 -696 579
rect -660 585 -648 588
rect -660 579 -657 585
rect -651 579 -648 585
rect -708 555 -705 561
rect -699 555 -696 561
rect -708 549 -696 555
rect -708 543 -705 549
rect -699 543 -696 549
rect -708 537 -696 543
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 528 -696 531
rect -684 561 -672 564
rect -684 555 -681 561
rect -675 555 -672 561
rect -684 549 -672 555
rect -684 543 -681 549
rect -675 543 -672 549
rect -684 537 -672 543
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 489 -672 531
rect -660 561 -648 579
rect -612 585 -600 588
rect -612 579 -609 585
rect -603 579 -600 585
rect -660 555 -657 561
rect -651 555 -648 561
rect -660 549 -648 555
rect -660 543 -657 549
rect -651 543 -648 549
rect -660 537 -648 543
rect -660 531 -657 537
rect -651 531 -648 537
rect -660 528 -648 531
rect -636 561 -624 564
rect -636 555 -633 561
rect -627 555 -624 561
rect -636 549 -624 555
rect -636 543 -633 549
rect -627 543 -624 549
rect -636 537 -624 543
rect -636 531 -633 537
rect -627 531 -624 537
rect -660 513 -648 516
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 504 -648 507
rect -684 483 -681 489
rect -675 483 -672 489
rect -708 441 -696 444
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 417 -696 435
rect -684 441 -672 483
rect -636 489 -624 531
rect -612 561 -600 579
rect -612 555 -609 561
rect -603 555 -600 561
rect -612 549 -600 555
rect -612 543 -609 549
rect -603 543 -600 549
rect -612 537 -600 543
rect -612 531 -609 537
rect -603 531 -600 537
rect -612 528 -600 531
rect -636 483 -633 489
rect -627 483 -624 489
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 432 -672 435
rect -660 441 -648 444
rect -660 435 -657 441
rect -651 435 -648 441
rect -708 411 -705 417
rect -699 411 -696 417
rect -708 405 -696 411
rect -708 399 -705 405
rect -699 399 -696 405
rect -660 417 -648 435
rect -636 441 -624 483
rect -636 435 -633 441
rect -627 435 -624 441
rect -636 432 -624 435
rect -612 441 -600 444
rect -612 435 -609 441
rect -603 435 -600 441
rect -660 411 -657 417
rect -651 411 -648 417
rect -660 405 -648 411
rect -708 393 -696 399
rect -708 387 -705 393
rect -699 387 -696 393
rect -708 381 -696 387
rect -708 375 -705 381
rect -699 375 -696 381
rect -708 372 -696 375
rect -684 393 -672 402
rect -660 399 -657 405
rect -651 399 -648 405
rect -612 417 -600 435
rect -612 411 -609 417
rect -603 411 -600 417
rect -612 405 -600 411
rect -660 396 -648 399
rect -684 387 -681 393
rect -675 387 -672 393
rect -684 384 -672 387
rect -636 393 -624 402
rect -636 387 -633 393
rect -627 387 -624 393
rect -636 384 -624 387
rect -684 381 -624 384
rect -684 375 -681 381
rect -675 375 -633 381
rect -627 375 -624 381
rect -684 372 -624 375
rect -612 399 -609 405
rect -603 399 -600 405
rect -612 393 -600 399
rect -612 387 -609 393
rect -603 387 -600 393
rect -612 381 -600 387
rect -612 375 -609 381
rect -603 375 -600 381
rect -612 372 -600 375
rect -684 357 -672 360
rect -684 351 -681 357
rect -675 351 -672 357
rect -684 348 -672 351
rect -708 333 -696 336
rect -708 327 -705 333
rect -699 327 -696 333
rect -708 324 -696 327
rect -708 309 -696 312
rect -708 303 -705 309
rect -699 303 -696 309
rect -708 213 -696 303
rect -708 207 -705 213
rect -699 207 -696 213
rect -708 165 -696 207
rect -708 159 -705 165
rect -699 159 -696 165
rect -708 117 -696 159
rect -708 111 -705 117
rect -699 111 -696 117
rect -708 69 -696 111
rect -708 63 -705 69
rect -699 63 -696 69
rect -708 -27 -696 63
rect -708 -33 -705 -27
rect -699 -33 -696 -27
rect -708 -75 -696 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -123 -696 -105
rect -660 -75 -648 372
rect -636 357 -624 360
rect -636 351 -633 357
rect -627 351 -624 357
rect -636 348 -624 351
rect -612 333 -600 336
rect -612 327 -609 333
rect -603 327 -600 333
rect -612 324 -600 327
rect -612 309 -600 312
rect -612 303 -609 309
rect -603 303 -600 309
rect -612 213 -600 303
rect -612 207 -609 213
rect -603 207 -600 213
rect -612 165 -600 207
rect -612 159 -609 165
rect -603 159 -600 165
rect -612 117 -600 159
rect -612 111 -609 117
rect -603 111 -600 117
rect -612 69 -600 111
rect -612 63 -609 69
rect -603 63 -600 69
rect -612 -27 -600 63
rect -612 -33 -609 -27
rect -603 -33 -600 -27
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -612 -75 -600 -33
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -708 -129 -705 -123
rect -699 -129 -696 -123
rect -708 -132 -696 -129
rect -612 -123 -600 -105
rect -612 -129 -609 -123
rect -603 -129 -600 -123
rect -612 -132 -600 -129
<< via2 >>
rect -705 579 -699 585
rect -657 579 -651 585
rect -705 555 -699 561
rect -705 543 -699 549
rect -705 531 -699 537
rect -609 579 -603 585
rect -657 555 -651 561
rect -657 543 -651 549
rect -657 531 -651 537
rect -657 507 -651 513
rect -681 483 -675 489
rect -705 435 -699 441
rect -609 555 -603 561
rect -609 543 -603 549
rect -609 531 -603 537
rect -633 483 -627 489
rect -681 435 -675 441
rect -657 435 -651 441
rect -633 435 -627 441
rect -609 435 -603 441
rect -681 351 -675 357
rect -705 327 -699 333
rect -705 303 -699 309
rect -705 207 -699 213
rect -705 159 -699 165
rect -705 111 -699 117
rect -705 63 -699 69
rect -705 -33 -699 -27
rect -681 -57 -675 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -633 351 -627 357
rect -609 327 -603 333
rect -609 303 -603 309
rect -609 207 -603 213
rect -609 159 -603 165
rect -609 111 -603 117
rect -609 63 -603 69
rect -609 -33 -603 -27
rect -633 -57 -627 -51
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal3 >>
rect -720 585 -588 588
rect -720 579 -705 585
rect -699 579 -657 585
rect -651 579 -609 585
rect -603 579 -588 585
rect -720 561 -588 579
rect -720 555 -705 561
rect -699 555 -657 561
rect -651 555 -609 561
rect -603 555 -588 561
rect -720 549 -588 555
rect -720 543 -705 549
rect -699 543 -657 549
rect -651 543 -609 549
rect -603 543 -588 549
rect -720 537 -588 543
rect -720 531 -705 537
rect -699 531 -657 537
rect -651 531 -609 537
rect -603 531 -588 537
rect -720 528 -588 531
rect -660 513 -648 516
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 504 -648 507
rect -720 489 -588 492
rect -720 483 -681 489
rect -675 483 -633 489
rect -627 483 -588 489
rect -720 474 -588 483
rect -720 465 -588 468
rect -720 459 -657 465
rect -651 459 -588 465
rect -720 456 -588 459
rect -720 441 -588 450
rect -720 435 -705 441
rect -699 435 -681 441
rect -675 435 -657 441
rect -651 435 -633 441
rect -627 435 -609 441
rect -603 435 -588 441
rect -720 432 -588 435
rect -684 357 -672 360
rect -684 351 -681 357
rect -675 351 -672 357
rect -684 348 -672 351
rect -636 357 -624 360
rect -636 351 -633 357
rect -627 351 -624 357
rect -636 348 -624 351
rect -720 333 -588 336
rect -720 327 -705 333
rect -699 327 -609 333
rect -603 327 -588 333
rect -720 324 -588 327
rect -720 309 -588 312
rect -720 303 -705 309
rect -699 303 -609 309
rect -603 303 -588 309
rect -720 300 -588 303
rect -720 228 -588 288
rect -720 213 -588 216
rect -720 207 -705 213
rect -699 207 -609 213
rect -603 207 -588 213
rect -720 204 -588 207
rect -720 180 -588 192
rect -720 165 -588 168
rect -720 159 -705 165
rect -699 159 -609 165
rect -603 159 -588 165
rect -720 156 -588 159
rect -720 132 -588 144
rect -720 117 -588 120
rect -720 111 -705 117
rect -699 111 -609 117
rect -603 111 -588 117
rect -720 108 -588 111
rect -720 84 -588 96
rect -720 69 -588 72
rect -720 63 -705 69
rect -699 63 -609 69
rect -603 63 -588 69
rect -720 60 -588 63
rect -720 -12 -588 48
rect -720 -27 -588 -24
rect -720 -33 -705 -27
rect -699 -33 -609 -27
rect -603 -33 -588 -27
rect -720 -36 -588 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -720 -75 -588 -72
rect -720 -81 -705 -75
rect -699 -81 -609 -75
rect -603 -81 -588 -75
rect -720 -87 -588 -81
rect -720 -93 -705 -87
rect -699 -93 -609 -87
rect -603 -93 -588 -87
rect -720 -99 -588 -93
rect -720 -105 -705 -99
rect -699 -105 -609 -99
rect -603 -105 -588 -99
rect -720 -123 -588 -105
rect -720 -129 -705 -123
rect -699 -129 -609 -123
rect -603 -129 -588 -123
rect -720 -132 -588 -129
<< via3 >>
rect -657 507 -651 513
rect -681 483 -675 489
rect -633 483 -627 489
rect -657 459 -651 465
rect -705 435 -699 441
rect -681 435 -675 441
rect -633 435 -627 441
rect -609 435 -603 441
rect -681 351 -675 357
rect -633 351 -627 357
rect -681 -57 -675 -51
rect -633 -57 -627 -51
<< metal4 >>
rect -660 513 -648 516
rect -660 507 -657 513
rect -651 507 -648 513
rect -684 489 -672 492
rect -684 483 -681 489
rect -675 483 -672 489
rect -708 441 -696 444
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 432 -696 435
rect -684 441 -672 483
rect -660 465 -648 507
rect -660 459 -657 465
rect -651 459 -648 465
rect -660 456 -648 459
rect -636 489 -624 492
rect -636 483 -633 489
rect -627 483 -624 489
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 432 -672 435
rect -636 441 -624 483
rect -636 435 -633 441
rect -627 435 -624 441
rect -636 432 -624 435
rect -612 441 -600 444
rect -612 435 -609 441
rect -603 435 -600 441
rect -612 432 -600 435
rect -684 357 -672 360
rect -684 351 -681 357
rect -675 351 -672 357
rect -684 336 -672 351
rect -708 324 -672 336
rect -684 -51 -672 324
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 357 -624 360
rect -636 351 -633 357
rect -627 351 -624 357
rect -636 336 -624 351
rect -636 324 -600 336
rect -636 -51 -624 324
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
<< labels >>
rlabel metal4 -684 -12 -672 240 0 inl
port 1 nsew
rlabel metal4 -636 -12 -624 240 0 inr
port 2 nsew
rlabel metal2 -660 -12 -648 240 0 out
port 3 nsew
rlabel metal3 -720 528 -588 588 0 vdd
port 4 nsew
rlabel metal3 -720 456 -588 468 0 gp
port 5 nsew
rlabel nwell -720 324 -588 336 0 bp
port 6 nsew
rlabel metal3 -720 474 -708 492 0 vreg
port 7 nsew
rlabel metal3 -720 228 -588 288 0 op
port 8 nsew
rlabel metal3 -720 180 -588 192 0 im
port 9 nsew
rlabel metal3 -720 84 -588 96 0 ip
port 10 nsew
rlabel metal3 -720 -12 -588 48 0 om
port 11 nsew
rlabel metal3 -720 -132 -588 -72 0 gnd
port 12 nsew
rlabel metal1 -684 -108 -672 -72 0 d1
rlabel metal1 -636 -108 -624 -72 0 d2
rlabel metal1 -720 600 -588 612 0 vss
rlabel metal1 -720 456 -588 468 0 vss
<< end >>
