* NGSPICE file created from nautanauta.ext - technology: gf180mcuC

.subckt nautanauta_cell inl inr out gp vreg op xm im ip xp om vdd gnd bp
X0 vreg inr out bp pmos_3p3 w=1.5u l=0.6u
X1 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X2 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X3 out inr vreg bp pmos_3p3 w=1.5u l=0.6u
X4 dr inr out gnd nmos_3p3 w=1.8u l=0.6u
X5 vreg inl out bp pmos_3p3 w=1.5u l=0.6u
X6 dl inl gnd gnd nmos_3p3 w=1.8u l=0.6u
X7 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X8 gnd inr dr gnd nmos_3p3 w=1.8u l=0.6u
X9 out inl dl gnd nmos_3p3 w=1.8u l=0.6u
X10 out inl vreg bp pmos_3p3 w=1.5u l=0.6u
X11 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
C0 out inl 0.17fF
C1 bp inr 0.32fF
C2 vdd gp 0.66fF
C3 op inl 0.20fF
C4 out op 0.12fF
C5 vdd vreg 1.41fF
C6 om inr 0.18fF
C7 bp vreg 0.92fF
C8 bp inl 0.32fF
C9 gp vreg 1.98fF
C10 inl inr 0.55fF
C11 out bp 0.15fF
C12 out inr 0.19fF
C13 op inr 0.20fF
C14 xm op 1.35fF
C15 om inl 0.18fF
C16 out om 0.12fF
C17 out vreg 0.78fF
C18 xp om 1.35fF
C19 out gnd 1.48fF
C20 inr gnd 2.23fF
C21 inl gnd 2.25fF
C22 vreg gnd 0.72fF
C23 gp gnd 1.56fF
C24 bp gnd 6.58fF
C25 vdd gnd 6.08fF
C26 dr gnd 0.18fF
C27 dl gnd 0.18fF
.ends

.subckt nautanauta_edge gp vreg im ip xm op xp om vdd gnd bp
X0 gnd lo lo gnd nmos_3p3 w=1.8u l=0.6u
X1 vdd hih hih vdd pmos_6p0 w=1.8u l=0.6u
X2 vreg hi hi bp pmos_3p3 w=1.5u l=0.6u
C0 vreg gp 1.01fF
C1 hi vreg 0.11fF
C2 vdd vreg 0.22fF
C3 om xp 0.98fF
C4 hih vdd 0.45fF
C5 hi bp 0.28fF
C6 xm op 0.98fF
C7 bp vreg 0.23fF
C8 vreg gnd 0.44fF
C9 bp gnd 4.35fF
C10 vdd gnd 4.01fF
C11 lo gnd 0.84fF
C12 hi gnd 0.46fF
C13 hih gnd 0.46fF
.ends

.subckt nautanauta ip im op om vdd gp bp vreg gnd
Xnautanauta_cell_0 im im xp gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_1 xp xm xp gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_2 xm xp xm gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_3 ip ip xm gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_5 ip xp om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_4 xm im op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_6 om op om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_7 op om op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_8 xp ip om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_20 xm im op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_30 ip xp om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_31 xm im op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_9 im xm op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_21 ip xp om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_10 xm im op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_22 om op om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_11 ip xp om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_23 op om op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_12 om op om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_24 xp ip om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_13 op om op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_25 im xm op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_14 xp ip om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_26 im xm op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_15 im xm op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_16 im im xp gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_27 xp ip om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_17 xp xm xp gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_18 xm xp xm gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_28 op om op gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_29 om op om gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_cell_19 ip ip xm gp vreg op xm im ip xp om vdd gnd bp nautanauta_cell
Xnautanauta_edge_0 gp vreg im ip xm op xp om vdd gnd bp nautanauta_edge
Xnautanauta_edge_1 gp vreg im ip xm op xp om vdd gnd bp nautanauta_edge
X0 op xm mim_2p0fF c_width=199.2u c_length=7.2u
X1 om xp mim_2p0fF c_width=199.2u c_length=7.2u
C0 xm im 0.18fF
C1 vreg op 0.92fF
C2 op gp 0.50fF
C3 op om 1.03fF
C4 xm ip 1.22fF
C5 xm vdd 4.41fF
C6 om im 1.05fF
C7 op bp 0.15fF
C8 op xp 1.09fF
C9 vreg vdd 0.76fF
C10 vreg xm 0.82fF
C11 xp im 1.39fF
C12 om ip 0.93fF
C13 gp vdd 0.33fF
C14 xm gp 0.47fF
C15 om xm 0.80fF
C16 xp ip 0.87fF
C17 vreg gp -2.33fF
C18 vreg om 0.28fF
C19 op im 0.66fF
C20 xp xm 0.59fF
C21 vreg xp 0.15fF
C22 op ip 0.84fF
C23 op vdd 3.66fF
C24 ip im 3.03fF
C25 op xm 48.00fF
C26 xp om 50.34fF
C27 bp gnd 195.93fF
C28 im gnd 49.00fF
C29 vdd gnd 172.70fF
C30 om gnd 84.82fF
C31 ip gnd 48.71fF
C32 op gnd 69.88fF
C33 xm gnd 37.42fF
C34 xp gnd 42.15fF
C35 vreg gnd 8.66fF
C36 gp gnd 44.31fF
.ends

