* Amplifier open-loop DC testbench

* Include GF180MCU device models
.include "../../../gf180mcuC/libs.tech/ngspice/design.ngspice"
.lib "../../../gf180mcuC/libs.tech/ngspice/sm141064.ngspice" typical

.include "inv.spice"

.param pVDD = 5.0
.param pIB  = 20u

VDD vdd 0 dc {pVDD} pulse (0 {pVDD} 1n 100p 100p 1 1)
VSS vss 0 0
ECM cm vss vdd vss 0.5

ib vdd ib {pIB}
xb ib     vdd gp bp  vreg vss inv_bias
x0 in  out vdd gp bp  vreg vss inv0

.option gmin = 1e-15
.control

	dc vdd 1.0 6.0 10m
	plot vdd vreg gp vss xb.q ib
	plot xb.ref xb.q bp vreg
	
	wrdata ../data/inv_bias_vddsweep.txt vdd vreg gp
	
	dc ib 1u 100u 1u
	plot vreg
	
	tran 100p 40n uic
	plot vdd vreg gp
	wrdata ../data/inv_bias_tran.txt vdd vreg gp
.endc

.end
