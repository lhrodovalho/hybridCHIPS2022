magic
tech gf180mcuC
magscale 1 5
timestamp 1665184495
<< error_s >>
rect -5062 4202 -4598 4222
rect -5062 4194 -5042 4202
rect -5034 4194 -5006 4202
rect -4958 4194 -4930 4202
rect -4882 4194 -4854 4202
rect -4806 4194 -4778 4202
rect -4730 4194 -4702 4202
rect -4654 4194 -4626 4202
rect -4618 4194 -4598 4202
rect -5034 4166 -4986 4194
rect -4958 4166 -4910 4194
rect -4882 4166 -4834 4194
rect -4806 4166 -4758 4194
rect -4730 4166 -4682 4194
rect -4654 4166 -4598 4194
rect -5062 4118 -5042 4146
rect -5034 4118 -5006 4138
rect -4958 4118 -4930 4138
rect -4882 4118 -4854 4138
rect -4806 4118 -4778 4138
rect -4730 4118 -4702 4138
rect -4654 4118 -4626 4138
rect -4618 4118 -4598 4146
rect -5034 4090 -4986 4118
rect -4958 4090 -4910 4118
rect -4882 4090 -4834 4118
rect -4806 4090 -4758 4118
rect -4730 4090 -4682 4118
rect -4654 4090 -4598 4118
rect -5062 4042 -5042 4070
rect -5034 4042 -5006 4062
rect -4958 4042 -4930 4062
rect -4882 4042 -4854 4062
rect -4806 4042 -4778 4062
rect -4730 4042 -4702 4062
rect -4654 4042 -4626 4062
rect -4618 4042 -4598 4070
rect -5034 4014 -4986 4042
rect -4958 4014 -4910 4042
rect -4882 4014 -4834 4042
rect -4806 4014 -4758 4042
rect -4730 4014 -4682 4042
rect -4654 4014 -4598 4042
rect -5062 3966 -5042 3994
rect -5034 3966 -5006 3986
rect -4958 3966 -4930 3986
rect -4882 3966 -4854 3986
rect -4806 3966 -4778 3986
rect -4730 3966 -4702 3986
rect -4654 3966 -4626 3986
rect -4618 3966 -4598 3994
rect -5034 3938 -4986 3966
rect -4958 3938 -4910 3966
rect -4882 3938 -4834 3966
rect -4806 3938 -4758 3966
rect -4730 3938 -4682 3966
rect -4654 3938 -4598 3966
rect -5062 3890 -5042 3918
rect -5034 3890 -5006 3910
rect -4958 3890 -4930 3910
rect -4882 3890 -4854 3910
rect -4806 3890 -4778 3910
rect -4730 3890 -4702 3910
rect -4654 3890 -4626 3910
rect -4618 3890 -4598 3918
rect -5034 3862 -4986 3890
rect -4958 3862 -4910 3890
rect -4882 3862 -4834 3890
rect -4806 3862 -4758 3890
rect -4730 3862 -4682 3890
rect -4654 3862 -4598 3890
rect -5062 3814 -5042 3842
rect -5034 3814 -5006 3834
rect -4958 3814 -4930 3834
rect -4882 3814 -4854 3834
rect -4806 3814 -4778 3834
rect -4730 3814 -4702 3834
rect -4654 3814 -4626 3834
rect -4618 3814 -4598 3842
rect -5034 3786 -4986 3814
rect -4958 3786 -4910 3814
rect -4882 3786 -4834 3814
rect -4806 3786 -4758 3814
rect -4730 3786 -4682 3814
rect -4654 3786 -4598 3814
rect -5062 -1258 -4598 -1238
rect -5062 -1266 -5042 -1258
rect -5034 -1266 -5006 -1258
rect -4958 -1266 -4930 -1258
rect -4882 -1266 -4854 -1258
rect -4806 -1266 -4778 -1258
rect -4730 -1266 -4702 -1258
rect -4654 -1266 -4626 -1258
rect -4618 -1266 -4598 -1258
rect -5034 -1294 -4986 -1266
rect -4958 -1294 -4910 -1266
rect -4882 -1294 -4834 -1266
rect -4806 -1294 -4758 -1266
rect -4730 -1294 -4682 -1266
rect -4654 -1294 -4598 -1266
rect -5062 -1342 -5042 -1314
rect -5034 -1342 -5006 -1322
rect -4958 -1342 -4930 -1322
rect -4882 -1342 -4854 -1322
rect -4806 -1342 -4778 -1322
rect -4730 -1342 -4702 -1322
rect -4654 -1342 -4626 -1322
rect -4618 -1342 -4598 -1314
rect -5034 -1370 -4986 -1342
rect -4958 -1370 -4910 -1342
rect -4882 -1370 -4834 -1342
rect -4806 -1370 -4758 -1342
rect -4730 -1370 -4682 -1342
rect -4654 -1370 -4598 -1342
rect -5062 -1418 -5042 -1390
rect -5034 -1418 -5006 -1398
rect -4958 -1418 -4930 -1398
rect -4882 -1418 -4854 -1398
rect -4806 -1418 -4778 -1398
rect -4730 -1418 -4702 -1398
rect -4654 -1418 -4626 -1398
rect -4618 -1418 -4598 -1390
rect -5034 -1446 -4986 -1418
rect -4958 -1446 -4910 -1418
rect -4882 -1446 -4834 -1418
rect -4806 -1446 -4758 -1418
rect -4730 -1446 -4682 -1418
rect -4654 -1446 -4598 -1418
rect -5062 -1494 -5042 -1466
rect -5034 -1494 -5006 -1474
rect -4958 -1494 -4930 -1474
rect -4882 -1494 -4854 -1474
rect -4806 -1494 -4778 -1474
rect -4730 -1494 -4702 -1474
rect -4654 -1494 -4626 -1474
rect -4618 -1494 -4598 -1466
rect -5034 -1522 -4986 -1494
rect -4958 -1522 -4910 -1494
rect -4882 -1522 -4834 -1494
rect -4806 -1522 -4758 -1494
rect -4730 -1522 -4682 -1494
rect -4654 -1522 -4598 -1494
rect -5062 -1570 -5042 -1542
rect -5034 -1570 -5006 -1550
rect -4958 -1570 -4930 -1550
rect -4882 -1570 -4854 -1550
rect -4806 -1570 -4778 -1550
rect -4730 -1570 -4702 -1550
rect -4654 -1570 -4626 -1550
rect -4618 -1570 -4598 -1542
rect -5034 -1598 -4986 -1570
rect -4958 -1598 -4910 -1570
rect -4882 -1598 -4834 -1570
rect -4806 -1598 -4758 -1570
rect -4730 -1598 -4682 -1570
rect -4654 -1598 -4598 -1570
rect -5062 -1646 -5042 -1618
rect -5034 -1646 -5006 -1626
rect -4958 -1646 -4930 -1626
rect -4882 -1646 -4854 -1626
rect -4806 -1646 -4778 -1626
rect -4730 -1646 -4702 -1626
rect -4654 -1646 -4626 -1626
rect -4618 -1646 -4598 -1618
rect -5034 -1674 -4986 -1646
rect -4958 -1674 -4910 -1646
rect -4882 -1674 -4834 -1646
rect -4806 -1674 -4758 -1646
rect -4730 -1674 -4682 -1646
rect -4654 -1674 -4598 -1646
<< metal2 >>
rect -3840 1720 -3780 1740
rect -3840 1640 -3824 1720
rect -3796 1640 -3780 1720
rect -3840 1620 -3780 1640
rect -3240 1720 -3180 1740
rect -3240 1640 -3224 1720
rect -3196 1640 -3180 1720
rect -3240 1620 -3180 1640
rect 3960 1720 4020 1740
rect 3960 1640 3976 1720
rect 4004 1640 4020 1720
rect 3960 1620 4020 1640
rect 4560 1720 4620 1740
rect 4560 1640 4576 1720
rect 4604 1640 4620 1720
rect 4560 1620 4620 1640
rect 6360 1720 6420 1740
rect 6360 1640 6376 1720
rect 6404 1640 6420 1720
rect 6360 1620 6420 1640
rect 6960 1720 7020 1740
rect 6960 1640 6976 1720
rect 7004 1640 7020 1720
rect 6960 1620 7020 1640
rect 14160 1720 14220 1740
rect 14160 1640 14176 1720
rect 14204 1640 14220 1720
rect 14160 1620 14220 1640
rect 14760 1720 14820 1740
rect 14760 1640 14776 1720
rect 14804 1640 14820 1720
rect 14760 1620 14820 1640
rect -1440 1544 -1380 1560
rect -1440 1516 -1424 1544
rect -1396 1516 -1380 1544
rect -1440 1500 -1380 1516
rect 2160 1544 2220 1560
rect 2160 1516 2176 1544
rect 2204 1516 2220 1544
rect 2160 1500 2220 1516
rect 8760 1544 8820 1560
rect 8760 1516 8776 1544
rect 8804 1516 8820 1544
rect 8760 1500 8820 1516
rect 12360 1544 12420 1560
rect 12360 1516 12376 1544
rect 12404 1516 12420 1544
rect 12360 1500 12420 1516
rect -3840 1420 -3780 1440
rect -3840 1340 -3824 1420
rect -3796 1340 -3780 1420
rect -3840 1320 -3780 1340
rect -3240 1420 -3180 1440
rect -3240 1340 -3224 1420
rect -3196 1340 -3180 1420
rect -3240 1320 -3180 1340
rect 3960 1420 4020 1440
rect 3960 1340 3976 1420
rect 4004 1340 4020 1420
rect 3960 1320 4020 1340
rect 4560 1420 4620 1440
rect 4560 1340 4576 1420
rect 4604 1340 4620 1420
rect 4560 1320 4620 1340
rect 6360 1420 6420 1440
rect 6360 1340 6376 1420
rect 6404 1340 6420 1420
rect 6360 1320 6420 1340
rect 6960 1420 7020 1440
rect 6960 1340 6976 1420
rect 7004 1340 7020 1420
rect 6960 1320 7020 1340
rect 14160 1420 14220 1440
rect 14160 1340 14176 1420
rect 14204 1340 14220 1420
rect 14160 1320 14220 1340
rect 14760 1420 14820 1440
rect 14760 1340 14776 1420
rect 14804 1340 14820 1420
rect 14760 1320 14820 1340
rect -840 884 -780 900
rect -840 856 -824 884
rect -796 856 -780 884
rect -840 840 -780 856
rect 1560 884 1620 900
rect 1560 856 1576 884
rect 1604 856 1620 884
rect 1560 840 1620 856
rect 9360 884 9420 900
rect 9360 856 9376 884
rect 9404 856 9420 884
rect 9360 840 9420 856
rect 11760 884 11820 900
rect 11760 856 11776 884
rect 11804 856 11820 884
rect 11760 840 11820 856
rect -240 644 -180 660
rect -240 616 -224 644
rect -196 616 -180 644
rect -240 600 -180 616
rect 360 644 420 660
rect 360 616 376 644
rect 404 616 420 644
rect 360 600 420 616
rect 960 644 1020 660
rect 960 616 976 644
rect 1004 616 1020 644
rect 960 600 1020 616
rect 9960 644 10020 660
rect 9960 616 9976 644
rect 10004 616 10020 644
rect 9960 600 10020 616
rect 10560 644 10620 660
rect 10560 616 10576 644
rect 10604 616 10620 644
rect 10560 600 10620 616
rect 11160 644 11220 660
rect 11160 616 11176 644
rect 11204 616 11220 644
rect 11160 600 11220 616
rect -4440 160 -4380 180
rect -4440 80 -4424 160
rect -4396 80 -4380 160
rect -4440 60 -4380 80
rect -2640 160 -2580 180
rect -2640 80 -2624 160
rect -2596 80 -2580 160
rect -2640 60 -2580 80
rect 3360 160 3420 180
rect 3360 80 3376 160
rect 3404 80 3420 160
rect 3360 60 3420 80
rect 5160 160 5220 180
rect 5160 80 5176 160
rect 5204 80 5220 160
rect 5160 60 5220 80
rect 5760 160 5820 180
rect 5760 80 5776 160
rect 5804 80 5820 160
rect 5760 60 5820 80
rect 7560 160 7620 180
rect 7560 80 7576 160
rect 7604 80 7620 160
rect 7560 60 7620 80
rect 13560 160 13620 180
rect 13560 80 13576 160
rect 13604 80 13620 160
rect 13560 60 13620 80
rect 15360 160 15420 180
rect 15360 80 15376 160
rect 15404 80 15420 160
rect 15360 60 15420 80
rect -2040 -16 -1980 0
rect -2040 -44 -2024 -16
rect -1996 -44 -1980 -16
rect -2040 -60 -1980 -44
rect 2760 -16 2820 0
rect 2760 -44 2776 -16
rect 2804 -44 2820 -16
rect 2760 -60 2820 -44
rect 8160 -16 8220 0
rect 8160 -44 8176 -16
rect 8204 -44 8220 -16
rect 8160 -60 8220 -44
rect 12960 -16 13020 0
rect 12960 -44 12976 -16
rect 13004 -44 13020 -16
rect 12960 -60 13020 -44
rect -4440 -140 -4380 -120
rect -4440 -220 -4424 -140
rect -4396 -220 -4380 -140
rect -4440 -240 -4380 -220
rect -2640 -140 -2580 -120
rect -2640 -220 -2624 -140
rect -2596 -220 -2580 -140
rect -2640 -240 -2580 -220
rect 3360 -140 3420 -120
rect 3360 -220 3376 -140
rect 3404 -220 3420 -140
rect 3360 -240 3420 -220
rect 5160 -140 5220 -120
rect 5160 -220 5176 -140
rect 5204 -220 5220 -140
rect 5160 -240 5220 -220
rect 5760 -140 5820 -120
rect 5760 -220 5776 -140
rect 5804 -220 5820 -140
rect 5760 -240 5820 -220
rect 7560 -140 7620 -120
rect 7560 -220 7576 -140
rect 7604 -220 7620 -140
rect 7560 -240 7620 -220
rect 13560 -140 13620 -120
rect 13560 -220 13576 -140
rect 13604 -220 13620 -140
rect 13560 -240 13620 -220
rect 15360 -140 15420 -120
rect 15360 -220 15376 -140
rect 15404 -220 15420 -140
rect 15360 -240 15420 -220
<< via2 >>
rect -3824 1640 -3796 1720
rect -3224 1640 -3196 1720
rect 3976 1640 4004 1720
rect 4576 1640 4604 1720
rect 6376 1640 6404 1720
rect 6976 1640 7004 1720
rect 14176 1640 14204 1720
rect 14776 1640 14804 1720
rect -1424 1516 -1396 1544
rect 2176 1516 2204 1544
rect 8776 1516 8804 1544
rect 12376 1516 12404 1544
rect -3824 1340 -3796 1420
rect -3224 1340 -3196 1420
rect 3976 1340 4004 1420
rect 4576 1340 4604 1420
rect 6376 1340 6404 1420
rect 6976 1340 7004 1420
rect 14176 1340 14204 1420
rect 14776 1340 14804 1420
rect -824 856 -796 884
rect 1576 856 1604 884
rect 9376 856 9404 884
rect 11776 856 11804 884
rect -224 616 -196 644
rect 376 616 404 644
rect 976 616 1004 644
rect 9976 616 10004 644
rect 10576 616 10604 644
rect 11176 616 11204 644
rect -4424 80 -4396 160
rect -2624 80 -2596 160
rect 3376 80 3404 160
rect 5176 80 5204 160
rect 5776 80 5804 160
rect 7576 80 7604 160
rect 13576 80 13604 160
rect 15376 80 15404 160
rect -2024 -44 -1996 -16
rect 2776 -44 2804 -16
rect 8176 -44 8204 -16
rect 12976 -44 13004 -16
rect -4424 -220 -4396 -140
rect -2624 -220 -2596 -140
rect 3376 -220 3404 -140
rect 5176 -220 5204 -140
rect 5776 -220 5804 -140
rect 7576 -220 7604 -140
rect 13576 -220 13604 -140
rect 15376 -220 15404 -140
<< mimcap >>
rect -5100 4202 14880 4440
rect -5100 3778 -5042 4202
rect -4618 3778 14880 4202
rect -5100 3720 14880 3778
rect -5100 -1258 14880 -1200
rect -5100 -1682 -5042 -1258
rect -4618 -1682 14880 -1258
rect -5100 -1920 14880 -1682
<< mimcapcontact >>
rect -5042 3778 -4618 4202
rect -5042 -1682 -4618 -1258
<< metal3 >>
rect -5220 2940 -5160 3240
rect -5220 2670 -5160 2760
rect -5220 2580 -5160 2640
rect -5220 1920 -5160 1980
rect -5520 1705 -5160 1740
rect -5520 1625 -5504 1705
rect -5476 1625 -5264 1705
rect -5236 1625 -5160 1705
rect -5520 1590 -5160 1625
rect -3840 1720 -3780 1740
rect -3840 1640 -3824 1720
rect -3796 1640 -3780 1720
rect -3840 1620 -3780 1640
rect -3240 1720 -3180 1740
rect -3240 1640 -3224 1720
rect -3196 1640 -3180 1720
rect -3240 1620 -3180 1640
rect 840 1720 900 1740
rect 840 1640 856 1720
rect 884 1640 900 1720
rect 840 1620 900 1640
rect 3960 1720 4020 1740
rect 3960 1640 3976 1720
rect 4004 1640 4020 1720
rect 3960 1620 4020 1640
rect 4560 1720 4620 1740
rect 4560 1640 4576 1720
rect 4604 1640 4620 1720
rect 4560 1620 4620 1640
rect 6360 1720 6420 1740
rect 6360 1640 6376 1720
rect 6404 1640 6420 1720
rect 6360 1620 6420 1640
rect 6960 1720 7020 1740
rect 6960 1640 6976 1720
rect 7004 1640 7020 1720
rect 6960 1620 7020 1640
rect 10080 1720 10140 1740
rect 10080 1640 10096 1720
rect 10124 1640 10140 1720
rect 10080 1620 10140 1640
rect 14160 1720 14220 1740
rect 14160 1640 14176 1720
rect 14204 1640 14220 1720
rect 14160 1620 14220 1640
rect 14760 1720 14820 1740
rect 14760 1640 14776 1720
rect 14804 1640 14820 1720
rect 14760 1620 14820 1640
rect -5520 1544 -5160 1560
rect -5520 1516 -5384 1544
rect -5356 1516 -5160 1544
rect -5520 1500 -5160 1516
rect -3720 1544 -3660 1560
rect -3720 1516 -3704 1544
rect -3676 1516 -3660 1544
rect -3720 1500 -3660 1516
rect -3360 1544 -3300 1560
rect -3360 1516 -3344 1544
rect -3316 1516 -3300 1544
rect -3360 1500 -3300 1516
rect -1440 1544 -1380 1560
rect -1440 1516 -1424 1544
rect -1396 1516 -1380 1544
rect -1440 1500 -1380 1516
rect 1680 1544 1740 1560
rect 1680 1516 1696 1544
rect 1724 1516 1740 1544
rect 1680 1500 1740 1516
rect 2160 1544 2220 1560
rect 2160 1516 2176 1544
rect 2204 1516 2220 1544
rect 2160 1500 2220 1516
rect 4080 1544 4140 1560
rect 4080 1516 4096 1544
rect 4124 1516 4140 1544
rect 4080 1500 4140 1516
rect 4440 1544 4500 1560
rect 4440 1516 4456 1544
rect 4484 1516 4500 1544
rect 4440 1500 4500 1516
rect 6480 1544 6540 1560
rect 6480 1516 6496 1544
rect 6524 1516 6540 1544
rect 6480 1500 6540 1516
rect 6840 1544 6900 1560
rect 6840 1516 6856 1544
rect 6884 1516 6900 1544
rect 6840 1500 6900 1516
rect 8760 1544 8820 1560
rect 8760 1516 8776 1544
rect 8804 1516 8820 1544
rect 8760 1500 8820 1516
rect 9240 1544 9300 1560
rect 9240 1516 9256 1544
rect 9284 1516 9300 1544
rect 9240 1500 9300 1516
rect 12360 1544 12420 1560
rect 12360 1516 12376 1544
rect 12404 1516 12420 1544
rect 12360 1500 12420 1516
rect 14280 1544 14340 1560
rect 14280 1516 14296 1544
rect 14324 1516 14340 1544
rect 14280 1500 14340 1516
rect 14640 1544 14700 1560
rect 14640 1516 14656 1544
rect 14684 1516 14700 1544
rect 14640 1500 14700 1516
rect -5520 1435 -5160 1470
rect -5520 1355 -5504 1435
rect -5476 1355 -5264 1435
rect -5236 1355 -5160 1435
rect -5520 1320 -5160 1355
rect -3840 1420 -3780 1440
rect -3840 1340 -3824 1420
rect -3796 1340 -3780 1420
rect -3840 1320 -3780 1340
rect -3240 1420 -3180 1440
rect -3240 1340 -3224 1420
rect -3196 1340 -3180 1420
rect -3240 1320 -3180 1340
rect 840 1420 900 1440
rect 840 1340 856 1420
rect 884 1340 900 1420
rect 840 1320 900 1340
rect 3960 1420 4020 1440
rect 3960 1340 3976 1420
rect 4004 1340 4020 1420
rect 3960 1320 4020 1340
rect 4560 1420 4620 1440
rect 4560 1340 4576 1420
rect 4604 1340 4620 1420
rect 4560 1320 4620 1340
rect 6360 1420 6420 1440
rect 6360 1340 6376 1420
rect 6404 1340 6420 1420
rect 6360 1320 6420 1340
rect 6960 1420 7020 1440
rect 6960 1340 6976 1420
rect 7004 1340 7020 1420
rect 6960 1320 7020 1340
rect 10080 1420 10140 1440
rect 10080 1340 10096 1420
rect 10124 1340 10140 1420
rect 10080 1320 10140 1340
rect 14160 1420 14220 1440
rect 14160 1340 14176 1420
rect 14204 1340 14220 1420
rect 14160 1320 14220 1340
rect 14760 1420 14820 1440
rect 14760 1340 14776 1420
rect 14804 1340 14820 1420
rect 14760 1320 14820 1340
rect -5220 1080 -5160 1140
rect -3960 1124 -3900 1140
rect -3960 1096 -3944 1124
rect -3916 1096 -3900 1124
rect -3960 1080 -3900 1096
rect -3120 1124 -3060 1140
rect -3120 1096 -3104 1124
rect -3076 1096 -3060 1124
rect -3120 1080 -3060 1096
rect -2160 1124 -2100 1140
rect -2160 1096 -2144 1124
rect -2116 1096 -2100 1124
rect -2160 1080 -2100 1096
rect 2880 1124 2940 1140
rect 2880 1096 2896 1124
rect 2924 1096 2940 1124
rect 2880 1080 2940 1096
rect 3840 1124 3900 1140
rect 3840 1096 3856 1124
rect 3884 1096 3900 1124
rect 3840 1080 3900 1096
rect 4680 1124 4740 1140
rect 4680 1096 4696 1124
rect 4724 1096 4740 1124
rect 4680 1080 4740 1096
rect 6240 1124 6300 1140
rect 6240 1096 6256 1124
rect 6284 1096 6300 1124
rect 6240 1080 6300 1096
rect 7080 1124 7140 1140
rect 7080 1096 7096 1124
rect 7124 1096 7140 1124
rect 7080 1080 7140 1096
rect 8040 1124 8100 1140
rect 8040 1096 8056 1124
rect 8084 1096 8100 1124
rect 8040 1080 8100 1096
rect 13080 1124 13140 1140
rect 13080 1096 13096 1124
rect 13124 1096 13140 1124
rect 13080 1080 13140 1096
rect 14040 1124 14100 1140
rect 14040 1096 14056 1124
rect 14084 1096 14100 1124
rect 14040 1080 14100 1096
rect 14880 1124 14940 1140
rect 14880 1096 14896 1124
rect 14924 1096 14940 1124
rect 14880 1080 14940 1096
rect -5220 840 -5160 900
rect -840 884 -780 900
rect -840 856 -824 884
rect -796 856 -780 884
rect -840 840 -780 856
rect -720 884 -660 900
rect -720 856 -704 884
rect -676 856 -660 884
rect -720 840 -660 856
rect -360 884 -300 900
rect -360 856 -344 884
rect -316 856 -300 884
rect -360 840 -300 856
rect 1080 884 1140 900
rect 1080 856 1096 884
rect 1124 856 1140 884
rect 1080 840 1140 856
rect 1440 884 1500 900
rect 1440 856 1456 884
rect 1484 856 1500 884
rect 1440 840 1500 856
rect 1560 884 1620 900
rect 1560 856 1576 884
rect 1604 856 1620 884
rect 1560 840 1620 856
rect 9360 884 9420 900
rect 9360 856 9376 884
rect 9404 856 9420 884
rect 9360 840 9420 856
rect 9480 884 9540 900
rect 9480 856 9496 884
rect 9524 856 9540 884
rect 9480 840 9540 856
rect 9840 884 9900 900
rect 9840 856 9856 884
rect 9884 856 9900 884
rect 9840 840 9900 856
rect 11280 884 11340 900
rect 11280 856 11296 884
rect 11324 856 11340 884
rect 11280 840 11340 856
rect 11640 884 11700 900
rect 11640 856 11656 884
rect 11684 856 11700 884
rect 11640 840 11700 856
rect 11760 884 11820 900
rect 11760 856 11776 884
rect 11804 856 11820 884
rect 11760 840 11820 856
rect -5220 600 -5160 660
rect -1920 644 -1860 660
rect -1920 616 -1904 644
rect -1876 616 -1860 644
rect -1920 600 -1860 616
rect -1560 644 -1500 660
rect -1560 616 -1544 644
rect -1516 616 -1500 644
rect -1560 600 -1500 616
rect -240 644 -180 660
rect -240 616 -224 644
rect -196 616 -180 644
rect -240 600 -180 616
rect 240 644 300 660
rect 240 616 256 644
rect 284 616 300 644
rect 240 600 300 616
rect 360 644 420 660
rect 360 616 376 644
rect 404 616 420 644
rect 360 600 420 616
rect 480 644 540 660
rect 480 616 496 644
rect 524 616 540 644
rect 480 600 540 616
rect 960 644 1020 660
rect 960 616 976 644
rect 1004 616 1020 644
rect 960 600 1020 616
rect 2280 644 2340 660
rect 2280 616 2296 644
rect 2324 616 2340 644
rect 2280 600 2340 616
rect 2640 644 2700 660
rect 2640 616 2656 644
rect 2684 616 2700 644
rect 2640 600 2700 616
rect 8280 644 8340 660
rect 8280 616 8296 644
rect 8324 616 8340 644
rect 8280 600 8340 616
rect 8640 644 8700 660
rect 8640 616 8656 644
rect 8684 616 8700 644
rect 8640 600 8700 616
rect 9960 644 10020 660
rect 9960 616 9976 644
rect 10004 616 10020 644
rect 9960 600 10020 616
rect 10440 644 10500 660
rect 10440 616 10456 644
rect 10484 616 10500 644
rect 10440 600 10500 616
rect 10560 644 10620 660
rect 10560 616 10576 644
rect 10604 616 10620 644
rect 10560 600 10620 616
rect 10680 644 10740 660
rect 10680 616 10696 644
rect 10724 616 10740 644
rect 10680 600 10740 616
rect 11160 644 11220 660
rect 11160 616 11176 644
rect 11204 616 11220 644
rect 11160 600 11220 616
rect 12480 644 12540 660
rect 12480 616 12496 644
rect 12524 616 12540 644
rect 12480 600 12540 616
rect 12840 644 12900 660
rect 12840 616 12856 644
rect 12884 616 12900 644
rect 12840 600 12900 616
rect -5220 360 -5160 420
rect -4320 404 -4260 420
rect -4320 376 -4304 404
rect -4276 376 -4260 404
rect -4320 360 -4260 376
rect -2760 404 -2700 420
rect -2760 376 -2744 404
rect -2716 376 -2700 404
rect -2760 360 -2700 376
rect -1320 404 -1260 420
rect -1320 376 -1304 404
rect -1276 376 -1260 404
rect -1320 360 -1260 376
rect 2040 404 2100 420
rect 2040 376 2056 404
rect 2084 376 2100 404
rect 2040 360 2100 376
rect 3480 404 3540 420
rect 3480 376 3496 404
rect 3524 376 3540 404
rect 3480 360 3540 376
rect 5040 404 5100 420
rect 5040 376 5056 404
rect 5084 376 5100 404
rect 5040 360 5100 376
rect 5880 404 5940 420
rect 5880 376 5896 404
rect 5924 376 5940 404
rect 5880 360 5940 376
rect 7440 404 7500 420
rect 7440 376 7456 404
rect 7484 376 7500 404
rect 7440 360 7500 376
rect 8880 404 8940 420
rect 8880 376 8896 404
rect 8924 376 8940 404
rect 8880 360 8940 376
rect 12240 404 12300 420
rect 12240 376 12256 404
rect 12284 376 12300 404
rect 12240 360 12300 376
rect 13680 404 13740 420
rect 13680 376 13696 404
rect 13724 376 13740 404
rect 13680 360 13740 376
rect 15240 404 15300 420
rect 15240 376 15256 404
rect 15284 376 15300 404
rect 15240 360 15300 376
rect -5520 145 -5160 180
rect -5520 65 -5504 145
rect -5476 65 -5264 145
rect -5236 65 -5160 145
rect -5520 30 -5160 65
rect -4440 160 -4380 180
rect -4440 80 -4424 160
rect -4396 80 -4380 160
rect -4440 60 -4380 80
rect -2640 160 -2580 180
rect -2640 80 -2624 160
rect -2596 80 -2580 160
rect -2640 60 -2580 80
rect -120 160 -60 180
rect -120 80 -104 160
rect -76 80 -60 160
rect -120 60 -60 80
rect 3360 160 3420 180
rect 3360 80 3376 160
rect 3404 80 3420 160
rect 3360 60 3420 80
rect 5160 160 5220 180
rect 5160 80 5176 160
rect 5204 80 5220 160
rect 5160 60 5220 80
rect 5760 160 5820 180
rect 5760 80 5776 160
rect 5804 80 5820 160
rect 5760 60 5820 80
rect 7560 160 7620 180
rect 7560 80 7576 160
rect 7604 80 7620 160
rect 7560 60 7620 80
rect 11040 160 11100 180
rect 11040 80 11056 160
rect 11084 80 11100 160
rect 11040 60 11100 80
rect 13560 160 13620 180
rect 13560 80 13576 160
rect 13604 80 13620 160
rect 13560 60 13620 80
rect 15360 160 15420 180
rect 15360 80 15376 160
rect 15404 80 15420 160
rect 15360 60 15420 80
rect -5520 -16 -5160 0
rect -5520 -44 -5384 -16
rect -5356 -44 -5160 -16
rect -5520 -60 -5160 -44
rect -4560 -16 -4500 0
rect -4560 -44 -4544 -16
rect -4516 -44 -4500 -16
rect -4560 -60 -4500 -44
rect -2520 -16 -2460 0
rect -2520 -44 -2504 -16
rect -2476 -44 -2460 -16
rect -2520 -60 -2460 -44
rect -2040 -16 -1980 0
rect -2040 -44 -2024 -16
rect -1996 -44 -1980 -16
rect -2040 -60 -1980 -44
rect -960 -16 -900 0
rect -960 -44 -944 -16
rect -916 -44 -900 -16
rect -960 -60 -900 -44
rect 2760 -16 2820 0
rect 2760 -44 2776 -16
rect 2804 -44 2820 -16
rect 2760 -60 2820 -44
rect 3240 -16 3300 0
rect 3240 -44 3256 -16
rect 3284 -44 3300 -16
rect 3240 -60 3300 -44
rect 5280 -16 5340 0
rect 5280 -44 5296 -16
rect 5324 -44 5340 -16
rect 5280 -60 5340 -44
rect 5640 -16 5700 0
rect 5640 -44 5656 -16
rect 5684 -44 5700 -16
rect 5640 -60 5700 -44
rect 7680 -16 7740 0
rect 7680 -44 7696 -16
rect 7724 -44 7740 -16
rect 7680 -60 7740 -44
rect 8160 -16 8220 0
rect 8160 -44 8176 -16
rect 8204 -44 8220 -16
rect 8160 -60 8220 -44
rect 11880 -16 11940 0
rect 11880 -44 11896 -16
rect 11924 -44 11940 -16
rect 11880 -60 11940 -44
rect 12960 -16 13020 0
rect 12960 -44 12976 -16
rect 13004 -44 13020 -16
rect 12960 -60 13020 -44
rect 13440 -16 13500 0
rect 13440 -44 13456 -16
rect 13484 -44 13500 -16
rect 13440 -60 13500 -44
rect 15480 -16 15540 0
rect 15480 -44 15496 -16
rect 15524 -44 15540 -16
rect 15480 -60 15540 -44
rect -5520 -125 -5160 -90
rect -5520 -205 -5504 -125
rect -5476 -205 -5264 -125
rect -5236 -205 -5160 -125
rect -5520 -240 -5160 -205
rect -4440 -140 -4380 -120
rect -4440 -220 -4424 -140
rect -4396 -220 -4380 -140
rect -4440 -240 -4380 -220
rect -2640 -140 -2580 -120
rect -2640 -220 -2624 -140
rect -2596 -220 -2580 -140
rect -2640 -240 -2580 -220
rect -120 -140 -60 -120
rect -120 -220 -104 -140
rect -76 -220 -60 -140
rect -120 -240 -60 -220
rect 3360 -140 3420 -120
rect 3360 -220 3376 -140
rect 3404 -220 3420 -140
rect 3360 -240 3420 -220
rect 5160 -140 5220 -120
rect 5160 -220 5176 -140
rect 5204 -220 5220 -140
rect 5160 -240 5220 -220
rect 5760 -140 5820 -120
rect 5760 -220 5776 -140
rect 5804 -220 5820 -140
rect 5760 -240 5820 -220
rect 7560 -140 7620 -120
rect 7560 -220 7576 -140
rect 7604 -220 7620 -140
rect 7560 -240 7620 -220
rect 11040 -140 11100 -120
rect 11040 -220 11056 -140
rect 11084 -220 11100 -140
rect 11040 -240 11100 -220
rect 13560 -140 13620 -120
rect 13560 -220 13576 -140
rect 13604 -220 13620 -140
rect 13560 -240 13620 -220
rect 15360 -140 15420 -120
rect 15360 -220 15376 -140
rect 15404 -220 15420 -140
rect 15360 -240 15420 -220
rect -5220 -840 -5160 -540
<< via3 >>
rect -5504 1625 -5476 1705
rect -5264 1625 -5236 1705
rect 856 1640 884 1720
rect 10096 1640 10124 1720
rect -5384 1516 -5356 1544
rect -3704 1516 -3676 1544
rect -3344 1516 -3316 1544
rect 1696 1516 1724 1544
rect 4096 1516 4124 1544
rect 4456 1516 4484 1544
rect 6496 1516 6524 1544
rect 6856 1516 6884 1544
rect 9256 1516 9284 1544
rect 14296 1516 14324 1544
rect 14656 1516 14684 1544
rect -5504 1355 -5476 1435
rect -5264 1355 -5236 1435
rect 856 1340 884 1420
rect 10096 1340 10124 1420
rect -3944 1096 -3916 1124
rect -3104 1096 -3076 1124
rect -2144 1096 -2116 1124
rect 2896 1096 2924 1124
rect 3856 1096 3884 1124
rect 4696 1096 4724 1124
rect 6256 1096 6284 1124
rect 7096 1096 7124 1124
rect 8056 1096 8084 1124
rect 13096 1096 13124 1124
rect 14056 1096 14084 1124
rect 14896 1096 14924 1124
rect -704 856 -676 884
rect -344 856 -316 884
rect 1096 856 1124 884
rect 1456 856 1484 884
rect 9496 856 9524 884
rect 9856 856 9884 884
rect 11296 856 11324 884
rect 11656 856 11684 884
rect -1904 616 -1876 644
rect -1544 616 -1516 644
rect 256 616 284 644
rect 496 616 524 644
rect 2296 616 2324 644
rect 2656 616 2684 644
rect 8296 616 8324 644
rect 8656 616 8684 644
rect 10456 616 10484 644
rect 10696 616 10724 644
rect 12496 616 12524 644
rect 12856 616 12884 644
rect -4304 376 -4276 404
rect -2744 376 -2716 404
rect -1304 376 -1276 404
rect 2056 376 2084 404
rect 3496 376 3524 404
rect 5056 376 5084 404
rect 5896 376 5924 404
rect 7456 376 7484 404
rect 8896 376 8924 404
rect 12256 376 12284 404
rect 13696 376 13724 404
rect 15256 376 15284 404
rect -5504 65 -5476 145
rect -5264 65 -5236 145
rect -104 80 -76 160
rect 11056 80 11084 160
rect -5384 -44 -5356 -16
rect -4544 -44 -4516 -16
rect -2504 -44 -2476 -16
rect -944 -44 -916 -16
rect 3256 -44 3284 -16
rect 5296 -44 5324 -16
rect 5656 -44 5684 -16
rect 7696 -44 7724 -16
rect 11896 -44 11924 -16
rect 13456 -44 13484 -16
rect 15496 -44 15524 -16
rect -5504 -205 -5476 -125
rect -5264 -205 -5236 -125
rect -104 -220 -76 -140
rect 11056 -220 11084 -140
<< metal4 >>
rect -5160 4440 14940 4500
rect -5520 3704 -5460 3780
rect -5520 3676 -5504 3704
rect -5476 3676 -5460 3704
rect -5520 3464 -5460 3676
rect -5520 3436 -5504 3464
rect -5476 3436 -5460 3464
rect -5520 1705 -5460 3436
rect -5520 1625 -5504 1705
rect -5476 1625 -5460 1705
rect -5520 1435 -5460 1625
rect -5520 1355 -5504 1435
rect -5476 1355 -5460 1435
rect -5520 1320 -5460 1355
rect -5400 3584 -5340 3780
rect -5400 3556 -5384 3584
rect -5356 3556 -5340 3584
rect -5400 1544 -5340 3556
rect -5400 1516 -5384 1544
rect -5356 1516 -5340 1544
rect -5400 1320 -5340 1516
rect -5280 3704 -5220 3780
rect -5280 3676 -5264 3704
rect -5236 3676 -5220 3704
rect -5280 3464 -5220 3676
rect -5160 3720 -5100 4440
rect 14880 3720 14940 4440
rect -5160 3584 14940 3720
rect -5160 3556 -5082 3584
rect 14862 3556 14940 3584
rect -5160 3540 14940 3556
rect -5280 3436 -5264 3464
rect -5236 3436 -5220 3464
rect -5280 1705 -5220 3436
rect -5280 1625 -5264 1705
rect -5236 1625 -5220 1705
rect -5280 1435 -5220 1625
rect 840 1720 900 1740
rect 840 1640 856 1720
rect 884 1640 900 1720
rect 840 1620 900 1640
rect 10080 1720 10140 1740
rect 10080 1640 10096 1720
rect 10124 1640 10140 1720
rect 10080 1620 10140 1640
rect -3720 1544 -3660 1560
rect -3720 1516 -3704 1544
rect -3676 1516 -3660 1544
rect -3720 1500 -3660 1516
rect -3360 1544 -3300 1560
rect -3360 1516 -3344 1544
rect -3316 1516 -3300 1544
rect -3360 1500 -3300 1516
rect 1680 1544 1740 1560
rect 1680 1516 1696 1544
rect 1724 1516 1740 1544
rect 1680 1500 1740 1516
rect 4080 1544 4140 1560
rect 4080 1516 4096 1544
rect 4124 1516 4140 1544
rect 4080 1500 4140 1516
rect 4440 1544 4500 1560
rect 4440 1516 4456 1544
rect 4484 1516 4500 1544
rect 4440 1500 4500 1516
rect 6480 1544 6540 1560
rect 6480 1516 6496 1544
rect 6524 1516 6540 1544
rect 6480 1500 6540 1516
rect 6840 1544 6900 1560
rect 6840 1516 6856 1544
rect 6884 1516 6900 1544
rect 6840 1500 6900 1516
rect 9240 1544 9300 1560
rect 9240 1516 9256 1544
rect 9284 1516 9300 1544
rect 9240 1500 9300 1516
rect 14280 1544 14340 1560
rect 14280 1516 14296 1544
rect 14324 1516 14340 1544
rect 14280 1500 14340 1516
rect 14640 1544 14700 1560
rect 14640 1516 14656 1544
rect 14684 1516 14700 1544
rect 14640 1500 14700 1516
rect -5280 1355 -5264 1435
rect -5236 1355 -5220 1435
rect -5280 1320 -5220 1355
rect 840 1420 900 1440
rect 840 1340 856 1420
rect 884 1340 900 1420
rect 840 1320 900 1340
rect 10080 1420 10140 1440
rect 10080 1340 10096 1420
rect 10124 1340 10140 1420
rect 10080 1320 10140 1340
rect -3960 1124 -3900 1140
rect -3960 1096 -3944 1124
rect -3916 1096 -3900 1124
rect -3960 1080 -3900 1096
rect -3120 1124 -3060 1140
rect -3120 1096 -3104 1124
rect -3076 1096 -3060 1124
rect -3120 1080 -3060 1096
rect -2160 1124 -2100 1140
rect -2160 1096 -2144 1124
rect -2116 1096 -2100 1124
rect -2160 1080 -2100 1096
rect 2880 1124 2940 1140
rect 2880 1096 2896 1124
rect 2924 1096 2940 1124
rect 2880 1080 2940 1096
rect 3840 1124 3900 1140
rect 3840 1096 3856 1124
rect 3884 1096 3900 1124
rect 3840 1080 3900 1096
rect 4680 1124 4740 1140
rect 4680 1096 4696 1124
rect 4724 1096 4740 1124
rect 4680 1080 4740 1096
rect 6240 1124 6300 1140
rect 6240 1096 6256 1124
rect 6284 1096 6300 1124
rect 6240 1080 6300 1096
rect 7080 1124 7140 1140
rect 7080 1096 7096 1124
rect 7124 1096 7140 1124
rect 7080 1080 7140 1096
rect 8040 1124 8100 1140
rect 8040 1096 8056 1124
rect 8084 1096 8100 1124
rect 8040 1080 8100 1096
rect 13080 1124 13140 1140
rect 13080 1096 13096 1124
rect 13124 1096 13140 1124
rect 13080 1080 13140 1096
rect 14040 1124 14100 1140
rect 14040 1096 14056 1124
rect 14084 1096 14100 1124
rect 14040 1080 14100 1096
rect 14880 1124 14940 1140
rect 14880 1096 14896 1124
rect 14924 1096 14940 1124
rect 14880 1080 14940 1096
rect -720 884 -660 900
rect -720 856 -704 884
rect -676 856 -660 884
rect -720 840 -660 856
rect -360 884 -300 900
rect -360 856 -344 884
rect -316 856 -300 884
rect -360 840 -300 856
rect 1080 884 1140 900
rect 1080 856 1096 884
rect 1124 856 1140 884
rect 1080 840 1140 856
rect 1440 884 1500 900
rect 1440 856 1456 884
rect 1484 856 1500 884
rect 1440 840 1500 856
rect 9480 884 9540 900
rect 9480 856 9496 884
rect 9524 856 9540 884
rect 9480 840 9540 856
rect 9840 884 9900 900
rect 9840 856 9856 884
rect 9884 856 9900 884
rect 9840 840 9900 856
rect 11280 884 11340 900
rect 11280 856 11296 884
rect 11324 856 11340 884
rect 11280 840 11340 856
rect 11640 884 11700 900
rect 11640 856 11656 884
rect 11684 856 11700 884
rect 11640 840 11700 856
rect -1920 644 -1860 660
rect -1920 616 -1904 644
rect -1876 616 -1860 644
rect -1920 600 -1860 616
rect -1560 644 -1500 660
rect -1560 616 -1544 644
rect -1516 616 -1500 644
rect -1560 600 -1500 616
rect 240 644 300 660
rect 240 616 256 644
rect 284 616 300 644
rect 240 600 300 616
rect 480 644 540 660
rect 480 616 496 644
rect 524 616 540 644
rect 480 600 540 616
rect 2280 644 2340 660
rect 2280 616 2296 644
rect 2324 616 2340 644
rect 2280 600 2340 616
rect 2640 644 2700 660
rect 2640 616 2656 644
rect 2684 616 2700 644
rect 2640 600 2700 616
rect 8280 644 8340 660
rect 8280 616 8296 644
rect 8324 616 8340 644
rect 8280 600 8340 616
rect 8640 644 8700 660
rect 8640 616 8656 644
rect 8684 616 8700 644
rect 8640 600 8700 616
rect 10440 644 10500 660
rect 10440 616 10456 644
rect 10484 616 10500 644
rect 10440 600 10500 616
rect 10680 644 10740 660
rect 10680 616 10696 644
rect 10724 616 10740 644
rect 10680 600 10740 616
rect 12480 644 12540 660
rect 12480 616 12496 644
rect 12524 616 12540 644
rect 12480 600 12540 616
rect 12840 644 12900 660
rect 12840 616 12856 644
rect 12884 616 12900 644
rect 12840 600 12900 616
rect -4320 404 -4260 420
rect -4320 376 -4304 404
rect -4276 376 -4260 404
rect -4320 360 -4260 376
rect -2760 404 -2700 420
rect -2760 376 -2744 404
rect -2716 376 -2700 404
rect -2760 360 -2700 376
rect -1320 404 -1260 420
rect -1320 376 -1304 404
rect -1276 376 -1260 404
rect -1320 360 -1260 376
rect 2040 404 2100 420
rect 2040 376 2056 404
rect 2084 376 2100 404
rect 2040 360 2100 376
rect 3480 404 3540 420
rect 3480 376 3496 404
rect 3524 376 3540 404
rect 3480 360 3540 376
rect 5040 404 5100 420
rect 5040 376 5056 404
rect 5084 376 5100 404
rect 5040 360 5100 376
rect 5880 404 5940 420
rect 5880 376 5896 404
rect 5924 376 5940 404
rect 5880 360 5940 376
rect 7440 404 7500 420
rect 7440 376 7456 404
rect 7484 376 7500 404
rect 7440 360 7500 376
rect 8880 404 8940 420
rect 8880 376 8896 404
rect 8924 376 8940 404
rect 8880 360 8940 376
rect 12240 404 12300 420
rect 12240 376 12256 404
rect 12284 376 12300 404
rect 12240 360 12300 376
rect 13680 404 13740 420
rect 13680 376 13696 404
rect 13724 376 13740 404
rect 13680 360 13740 376
rect 15240 404 15300 420
rect 15240 376 15256 404
rect 15284 376 15300 404
rect 15240 360 15300 376
rect -5520 145 -5460 180
rect -5520 65 -5504 145
rect -5476 65 -5460 145
rect -5520 -125 -5460 65
rect -5520 -205 -5504 -125
rect -5476 -205 -5460 -125
rect -5520 -916 -5460 -205
rect -5520 -944 -5504 -916
rect -5476 -944 -5460 -916
rect -5520 -1156 -5460 -944
rect -5520 -1184 -5504 -1156
rect -5476 -1184 -5460 -1156
rect -5520 -1260 -5460 -1184
rect -5400 -16 -5340 180
rect -5400 -44 -5384 -16
rect -5356 -44 -5340 -16
rect -5400 -1036 -5340 -44
rect -5400 -1064 -5384 -1036
rect -5356 -1064 -5340 -1036
rect -5400 -1260 -5340 -1064
rect -5280 145 -5220 180
rect -5280 65 -5264 145
rect -5236 65 -5220 145
rect -5280 -125 -5220 65
rect -120 160 -60 180
rect -120 80 -104 160
rect -76 80 -60 160
rect -120 60 -60 80
rect 11040 160 11100 180
rect 11040 80 11056 160
rect 11084 80 11100 160
rect 11040 60 11100 80
rect -4560 -16 -4500 0
rect -4560 -44 -4544 -16
rect -4516 -44 -4500 -16
rect -4560 -60 -4500 -44
rect -2520 -16 -2460 0
rect -2520 -44 -2504 -16
rect -2476 -44 -2460 -16
rect -2520 -60 -2460 -44
rect -960 -16 -900 0
rect -960 -44 -944 -16
rect -916 -44 -900 -16
rect -960 -60 -900 -44
rect 3240 -16 3300 0
rect 3240 -44 3256 -16
rect 3284 -44 3300 -16
rect 3240 -60 3300 -44
rect 5280 -16 5340 0
rect 5280 -44 5296 -16
rect 5324 -44 5340 -16
rect 5280 -60 5340 -44
rect 5640 -16 5700 0
rect 5640 -44 5656 -16
rect 5684 -44 5700 -16
rect 5640 -60 5700 -44
rect 7680 -16 7740 0
rect 7680 -44 7696 -16
rect 7724 -44 7740 -16
rect 7680 -60 7740 -44
rect 11880 -16 11940 0
rect 11880 -44 11896 -16
rect 11924 -44 11940 -16
rect 11880 -60 11940 -44
rect 13440 -16 13500 0
rect 13440 -44 13456 -16
rect 13484 -44 13500 -16
rect 13440 -60 13500 -44
rect 15480 -16 15540 0
rect 15480 -44 15496 -16
rect 15524 -44 15540 -16
rect 15480 -60 15540 -44
rect -5280 -205 -5264 -125
rect -5236 -205 -5220 -125
rect -5280 -916 -5220 -205
rect -120 -140 -60 -120
rect -120 -220 -104 -140
rect -76 -220 -60 -140
rect -120 -240 -60 -220
rect 11040 -140 11100 -120
rect 11040 -220 11056 -140
rect 11084 -220 11100 -140
rect 11040 -240 11100 -220
rect -5280 -944 -5264 -916
rect -5236 -944 -5220 -916
rect -5280 -1156 -5220 -944
rect -5280 -1184 -5264 -1156
rect -5236 -1184 -5220 -1156
rect -5280 -1260 -5220 -1184
rect -5160 -1036 14940 -1020
rect -5160 -1064 -5082 -1036
rect 14862 -1064 14940 -1036
rect -5160 -1200 14940 -1064
rect -5160 -1920 -5100 -1200
rect 14880 -1920 14940 -1200
rect -5160 -1980 14940 -1920
<< via4 >>
rect -5504 3676 -5476 3704
rect -5504 3436 -5476 3464
rect -5384 3556 -5356 3584
rect -5264 3676 -5236 3704
rect -5082 3556 14862 3584
rect -5264 3436 -5236 3464
rect -5504 -944 -5476 -916
rect -5504 -1184 -5476 -1156
rect -5384 -1064 -5356 -1036
rect -5264 -944 -5236 -916
rect -5264 -1184 -5236 -1156
rect -5082 -1064 14862 -1036
<< metal5 >>
rect -5160 4202 14940 4500
rect -5160 3778 -5042 4202
rect -5034 4166 -5006 4194
rect -4958 4166 -4930 4194
rect -4882 4166 -4854 4194
rect -4806 4166 -4778 4194
rect -4730 4166 -4702 4194
rect -4654 4166 -4626 4194
rect -5034 4090 -5006 4118
rect -4958 4090 -4930 4118
rect -4882 4090 -4854 4118
rect -4806 4090 -4778 4118
rect -4730 4090 -4702 4118
rect -4654 4090 -4626 4118
rect -5034 4014 -5006 4042
rect -4958 4014 -4930 4042
rect -4882 4014 -4854 4042
rect -4806 4014 -4778 4042
rect -4730 4014 -4702 4042
rect -4654 4014 -4626 4042
rect -5034 3938 -5006 3966
rect -4958 3938 -4930 3966
rect -4882 3938 -4854 3966
rect -4806 3938 -4778 3966
rect -4730 3938 -4702 3966
rect -4654 3938 -4626 3966
rect -5034 3862 -5006 3890
rect -4958 3862 -4930 3890
rect -4882 3862 -4854 3890
rect -4806 3862 -4778 3890
rect -4730 3862 -4702 3890
rect -4654 3862 -4626 3890
rect -5034 3786 -5006 3814
rect -4958 3786 -4930 3814
rect -4882 3786 -4854 3814
rect -4806 3786 -4778 3814
rect -4730 3786 -4702 3814
rect -4654 3786 -4626 3814
rect -4618 3778 14940 4202
rect -5160 3720 14940 3778
rect -5580 3704 14940 3720
rect -5580 3676 -5504 3704
rect -5476 3676 -5264 3704
rect -5236 3676 14940 3704
rect -5580 3660 14940 3676
rect -5580 3584 14940 3600
rect -5580 3556 -5384 3584
rect -5356 3556 -5082 3584
rect 14862 3556 14940 3584
rect -5580 3540 14940 3556
rect -5580 3464 14940 3480
rect -5580 3436 -5504 3464
rect -5476 3436 -5264 3464
rect -5236 3436 14940 3464
rect -5580 3420 14940 3436
rect -5580 -916 14940 -900
rect -5580 -944 -5504 -916
rect -5476 -944 -5264 -916
rect -5236 -944 14940 -916
rect -5580 -960 14940 -944
rect -5580 -1036 14940 -1020
rect -5580 -1064 -5384 -1036
rect -5356 -1064 -5082 -1036
rect 14862 -1064 14940 -1036
rect -5580 -1080 14940 -1064
rect -5580 -1156 14940 -1140
rect -5580 -1184 -5504 -1156
rect -5476 -1184 -5264 -1156
rect -5236 -1184 14940 -1156
rect -5580 -1200 14940 -1184
rect -5160 -1258 14940 -1200
rect -5160 -1682 -5042 -1258
rect -5034 -1294 -5006 -1266
rect -4958 -1294 -4930 -1266
rect -4882 -1294 -4854 -1266
rect -4806 -1294 -4778 -1266
rect -4730 -1294 -4702 -1266
rect -4654 -1294 -4626 -1266
rect -5034 -1370 -5006 -1342
rect -4958 -1370 -4930 -1342
rect -4882 -1370 -4854 -1342
rect -4806 -1370 -4778 -1342
rect -4730 -1370 -4702 -1342
rect -4654 -1370 -4626 -1342
rect -5034 -1446 -5006 -1418
rect -4958 -1446 -4930 -1418
rect -4882 -1446 -4854 -1418
rect -4806 -1446 -4778 -1418
rect -4730 -1446 -4702 -1418
rect -4654 -1446 -4626 -1418
rect -5034 -1522 -5006 -1494
rect -4958 -1522 -4930 -1494
rect -4882 -1522 -4854 -1494
rect -4806 -1522 -4778 -1494
rect -4730 -1522 -4702 -1494
rect -4654 -1522 -4626 -1494
rect -5034 -1598 -5006 -1570
rect -4958 -1598 -4930 -1570
rect -4882 -1598 -4854 -1570
rect -4806 -1598 -4778 -1570
rect -4730 -1598 -4702 -1570
rect -4654 -1598 -4626 -1570
rect -5034 -1674 -5006 -1646
rect -4958 -1674 -4930 -1646
rect -4882 -1674 -4854 -1646
rect -4806 -1674 -4778 -1646
rect -4730 -1674 -4702 -1646
rect -4654 -1674 -4626 -1646
rect -4618 -1682 14940 -1258
rect -5160 -1980 14940 -1682
use manfvieru_cell  manfvieru_cell_0
timestamp 1665184495
transform -1 0 12120 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_1
timestamp 1665184495
transform -1 0 11520 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_2
timestamp 1665184495
transform 1 0 17460 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_3
timestamp 1665184495
transform 1 0 16860 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_4
timestamp 1665184495
transform -1 0 9120 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_5
timestamp 1665184495
transform -1 0 9720 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_6
timestamp 1665184495
transform -1 0 8520 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_7
timestamp 1665184495
transform -1 0 7920 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_8
timestamp 1665184495
transform -1 0 7320 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_9
timestamp 1665184495
transform -1 0 6720 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_10
timestamp 1665184495
transform -1 0 6120 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_11
timestamp 1665184495
transform -1 0 5520 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_12
timestamp 1665184495
transform -1 0 4920 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_13
timestamp 1665184495
transform -1 0 4320 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_14
timestamp 1665184495
transform -1 0 3720 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_15
timestamp 1665184495
transform 1 0 9660 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_16
timestamp 1665184495
transform 1 0 9060 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_17
timestamp 1665184495
transform -1 0 1920 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_18
timestamp 1665184495
transform -1 0 1320 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_19
timestamp 1665184495
transform 1 0 7260 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_20
timestamp 1665184495
transform 1 0 6660 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_21
timestamp 1665184495
transform 1 0 6060 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_22
timestamp 1665184495
transform 1 0 5460 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_23
timestamp 1665184495
transform 1 0 4860 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_24
timestamp 1665184495
transform 1 0 4260 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_25
timestamp 1665184495
transform 1 0 3660 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_26
timestamp 1665184495
transform 1 0 3060 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_27
timestamp 1665184495
transform 1 0 2460 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_28
timestamp 1665184495
transform 1 0 1860 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_29
timestamp 1665184495
transform 1 0 1260 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_30
timestamp 1665184495
transform -1 0 -5880 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_31
timestamp 1665184495
transform -1 0 -6480 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_32
timestamp 1665184495
transform 1 0 -540 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_cell  manfvieru_cell_33
timestamp 1665184495
transform 1 0 -1140 0 1 -180
box -3600 -660 -2940 3540
use manfvieru_edge  manfvieru_edge_0
timestamp 1665184495
transform -1 0 12360 0 1 -180
box -3780 -660 -3300 3540
use manfvieru_edge  manfvieru_edge_1
timestamp 1665184495
transform 1 0 -1380 0 1 -180
box -3780 -660 -3300 3540
<< labels >>
rlabel metal3 s -5190 -30 -5190 -30 4 xp
rlabel metal3 s -5190 1530 -5190 1530 4 xm
rlabel metal3 s -5190 870 -5190 870 4 x
rlabel metal3 s -5190 630 -5190 630 4 y
rlabel metal3 s -5220 360 -5160 420 4 ip
port 1 nsew
rlabel metal3 s -5220 1080 -5160 1140 4 im
port 2 nsew
rlabel metal3 s -5220 1680 -5160 1740 4 op
port 3 nsew
rlabel metal3 s -5220 -240 -5160 -180 4 om
port 4 nsew
rlabel metal3 s -5220 2940 -5160 3240 4 vdd
port 5 nsew
rlabel metal3 s -5220 2580 -5160 2640 4 gp
port 6 nsew
rlabel metal3 s -5220 1920 -5160 1980 4 bp
port 7 nsew
rlabel metal3 s -5220 2700 -5160 2760 4 vreg
port 8 nsew
rlabel metal3 s -5220 -840 -5160 -540 4 gnd
port 9 nsew
<< end >>
