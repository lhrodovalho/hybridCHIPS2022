magic
tech gf180mcuC
magscale 1 5
timestamp 1665184495
<< error_p >>
rect 24818 5642 25282 5662
rect 24818 5634 24838 5642
rect 24846 5634 24874 5642
rect 24922 5634 24950 5642
rect 24998 5634 25026 5642
rect 25074 5634 25102 5642
rect 25150 5634 25178 5642
rect 25226 5634 25254 5642
rect 25262 5634 25282 5642
rect 24846 5606 24894 5634
rect 24922 5606 24970 5634
rect 24998 5606 25046 5634
rect 25074 5606 25122 5634
rect 25150 5606 25198 5634
rect 25226 5606 25282 5634
rect 24818 5558 24838 5586
rect 24846 5558 24874 5578
rect 24922 5558 24950 5578
rect 24998 5558 25026 5578
rect 25074 5558 25102 5578
rect 25150 5558 25178 5578
rect 25226 5558 25254 5578
rect 25262 5558 25282 5586
rect 24846 5530 24894 5558
rect 24922 5530 24970 5558
rect 24998 5530 25046 5558
rect 25074 5530 25122 5558
rect 25150 5530 25198 5558
rect 25226 5530 25282 5558
rect 24818 5482 24838 5510
rect 24846 5482 24874 5502
rect 24922 5482 24950 5502
rect 24998 5482 25026 5502
rect 25074 5482 25102 5502
rect 25150 5482 25178 5502
rect 25226 5482 25254 5502
rect 25262 5482 25282 5510
rect 24846 5454 24894 5482
rect 24922 5454 24970 5482
rect 24998 5454 25046 5482
rect 25074 5454 25122 5482
rect 25150 5454 25198 5482
rect 25226 5454 25282 5482
rect 24818 5406 24838 5434
rect 24846 5406 24874 5426
rect 24922 5406 24950 5426
rect 24998 5406 25026 5426
rect 25074 5406 25102 5426
rect 25150 5406 25178 5426
rect 25226 5406 25254 5426
rect 25262 5406 25282 5434
rect 24846 5378 24894 5406
rect 24922 5378 24970 5406
rect 24998 5378 25046 5406
rect 25074 5378 25122 5406
rect 25150 5378 25198 5406
rect 25226 5378 25282 5406
rect 24818 5330 24838 5358
rect 24846 5330 24874 5350
rect 24922 5330 24950 5350
rect 24998 5330 25026 5350
rect 25074 5330 25102 5350
rect 25150 5330 25178 5350
rect 25226 5330 25254 5350
rect 25262 5330 25282 5358
rect 24846 5302 24894 5330
rect 24922 5302 24970 5330
rect 24998 5302 25046 5330
rect 25074 5302 25122 5330
rect 25150 5302 25198 5330
rect 25226 5302 25282 5330
rect 24818 5254 24838 5282
rect 24846 5254 24874 5274
rect 24922 5254 24950 5274
rect 24998 5254 25026 5274
rect 25074 5254 25102 5274
rect 25150 5254 25178 5274
rect 25226 5254 25254 5274
rect 25262 5254 25282 5282
rect 24846 5226 24894 5254
rect 24922 5226 24970 5254
rect 24998 5226 25046 5254
rect 25074 5226 25122 5254
rect 25150 5226 25198 5254
rect 25226 5226 25282 5254
rect 24818 602 25282 622
rect 24818 594 24838 602
rect 24846 594 24874 602
rect 24922 594 24950 602
rect 24998 594 25026 602
rect 25074 594 25102 602
rect 25150 594 25178 602
rect 25226 594 25254 602
rect 25262 594 25282 602
rect 24846 580 24894 594
rect 24922 580 24970 594
rect 24998 580 25046 594
rect 25074 580 25122 594
rect 25150 580 25198 594
rect 25226 580 25282 594
rect 24846 -7854 24894 -7840
rect 24922 -7854 24970 -7840
rect 24998 -7854 25046 -7840
rect 25074 -7854 25122 -7840
rect 25150 -7854 25198 -7840
rect 25226 -7854 25282 -7840
rect 24818 -12898 25282 -12878
rect 24818 -12906 24838 -12898
rect 24846 -12906 24874 -12898
rect 24922 -12906 24950 -12898
rect 24998 -12906 25026 -12898
rect 25074 -12906 25102 -12898
rect 25150 -12906 25178 -12898
rect 25226 -12906 25254 -12898
rect 25262 -12906 25282 -12898
rect 24846 -12934 24894 -12906
rect 24922 -12934 24970 -12906
rect 24998 -12934 25046 -12906
rect 25074 -12934 25122 -12906
rect 25150 -12934 25198 -12906
rect 25226 -12934 25282 -12906
rect 24818 -12982 24838 -12954
rect 24846 -12982 24874 -12962
rect 24922 -12982 24950 -12962
rect 24998 -12982 25026 -12962
rect 25074 -12982 25102 -12962
rect 25150 -12982 25178 -12962
rect 25226 -12982 25254 -12962
rect 25262 -12982 25282 -12954
rect 24846 -13010 24894 -12982
rect 24922 -13010 24970 -12982
rect 24998 -13010 25046 -12982
rect 25074 -13010 25122 -12982
rect 25150 -13010 25198 -12982
rect 25226 -13010 25282 -12982
rect 24818 -13058 24838 -13030
rect 24846 -13058 24874 -13038
rect 24922 -13058 24950 -13038
rect 24998 -13058 25026 -13038
rect 25074 -13058 25102 -13038
rect 25150 -13058 25178 -13038
rect 25226 -13058 25254 -13038
rect 25262 -13058 25282 -13030
rect 24846 -13086 24894 -13058
rect 24922 -13086 24970 -13058
rect 24998 -13086 25046 -13058
rect 25074 -13086 25122 -13058
rect 25150 -13086 25198 -13058
rect 25226 -13086 25282 -13058
rect 24818 -13134 24838 -13106
rect 24846 -13134 24874 -13114
rect 24922 -13134 24950 -13114
rect 24998 -13134 25026 -13114
rect 25074 -13134 25102 -13114
rect 25150 -13134 25178 -13114
rect 25226 -13134 25254 -13114
rect 25262 -13134 25282 -13106
rect 24846 -13162 24894 -13134
rect 24922 -13162 24970 -13134
rect 24998 -13162 25046 -13134
rect 25074 -13162 25122 -13134
rect 25150 -13162 25198 -13134
rect 25226 -13162 25282 -13134
rect 24818 -13210 24838 -13182
rect 24846 -13210 24874 -13190
rect 24922 -13210 24950 -13190
rect 24998 -13210 25026 -13190
rect 25074 -13210 25102 -13190
rect 25150 -13210 25178 -13190
rect 25226 -13210 25254 -13190
rect 25262 -13210 25282 -13182
rect 24846 -13238 24894 -13210
rect 24922 -13238 24970 -13210
rect 24998 -13238 25046 -13210
rect 25074 -13238 25122 -13210
rect 25150 -13238 25198 -13210
rect 25226 -13238 25282 -13210
rect 24818 -13286 24838 -13258
rect 24846 -13286 24874 -13266
rect 24922 -13286 24950 -13266
rect 24998 -13286 25026 -13266
rect 25074 -13286 25102 -13266
rect 25150 -13286 25178 -13266
rect 25226 -13286 25254 -13266
rect 25262 -13286 25282 -13258
rect 24846 -13314 24894 -13286
rect 24922 -13314 24970 -13286
rect 24998 -13314 25046 -13286
rect 25074 -13314 25122 -13286
rect 25150 -13314 25198 -13286
rect 25226 -13314 25282 -13286
<< error_s >>
rect 24846 566 24894 580
rect 24922 566 24970 580
rect 24998 566 25046 580
rect 25074 566 25122 580
rect 25150 566 25198 580
rect 25226 566 25282 580
rect 24818 518 24838 546
rect 24846 518 24874 538
rect 24922 518 24950 538
rect 24998 518 25026 538
rect 25074 518 25102 538
rect 25150 518 25178 538
rect 25226 518 25254 538
rect 25262 518 25282 546
rect 24846 490 24894 518
rect 24922 490 24970 518
rect 24998 490 25046 518
rect 25074 490 25122 518
rect 25150 490 25198 518
rect 25226 490 25282 518
rect 24818 442 24838 470
rect 24846 442 24874 462
rect 24922 442 24950 462
rect 24998 442 25026 462
rect 25074 442 25102 462
rect 25150 442 25178 462
rect 25226 442 25254 462
rect 25262 442 25282 470
rect 24846 414 24894 442
rect 24922 414 24970 442
rect 24998 414 25046 442
rect 25074 414 25122 442
rect 25150 414 25198 442
rect 25226 414 25282 442
rect 24818 366 24838 394
rect 24846 366 24874 386
rect 24922 366 24950 386
rect 24998 366 25026 386
rect 25074 366 25102 386
rect 25150 366 25178 386
rect 25226 366 25254 386
rect 25262 366 25282 394
rect 24846 338 24894 366
rect 24922 338 24970 366
rect 24998 338 25046 366
rect 25074 338 25122 366
rect 25150 338 25198 366
rect 25226 338 25282 366
rect 24818 290 24838 318
rect 24846 290 24874 310
rect 24922 290 24950 310
rect 24998 290 25026 310
rect 25074 290 25102 310
rect 25150 290 25178 310
rect 25226 290 25254 310
rect 25262 290 25282 318
rect 24846 262 24894 290
rect 24922 262 24970 290
rect 24998 262 25046 290
rect 25074 262 25122 290
rect 25150 262 25198 290
rect 25226 262 25282 290
rect 24818 214 24838 242
rect 24846 214 24874 234
rect 24922 214 24950 234
rect 24998 214 25026 234
rect 25074 214 25102 234
rect 25150 214 25178 234
rect 25226 214 25254 234
rect 25262 214 25282 242
rect 24846 186 24894 214
rect 24922 186 24970 214
rect 24998 186 25046 214
rect 25074 186 25122 214
rect 25150 186 25198 214
rect 25226 186 25282 214
rect 25058 -898 25522 -878
rect 25058 -906 25078 -898
rect 25086 -906 25114 -898
rect 25162 -906 25190 -898
rect 25238 -906 25266 -898
rect 25314 -906 25342 -898
rect 25390 -906 25418 -898
rect 25466 -906 25494 -898
rect 25502 -906 25522 -898
rect 25086 -934 25134 -906
rect 25162 -934 25210 -906
rect 25238 -934 25286 -906
rect 25314 -934 25362 -906
rect 25390 -934 25438 -906
rect 25466 -934 25522 -906
rect 25058 -982 25078 -954
rect 25086 -982 25114 -962
rect 25162 -982 25190 -962
rect 25238 -982 25266 -962
rect 25314 -982 25342 -962
rect 25390 -982 25418 -962
rect 25466 -982 25494 -962
rect 25502 -982 25522 -954
rect 25086 -1010 25134 -982
rect 25162 -1010 25210 -982
rect 25238 -1010 25286 -982
rect 25314 -1010 25362 -982
rect 25390 -1010 25438 -982
rect 25466 -1010 25522 -982
rect 25058 -1058 25078 -1030
rect 25086 -1058 25114 -1038
rect 25162 -1058 25190 -1038
rect 25238 -1058 25266 -1038
rect 25314 -1058 25342 -1038
rect 25390 -1058 25418 -1038
rect 25466 -1058 25494 -1038
rect 25502 -1058 25522 -1030
rect 25086 -1086 25134 -1058
rect 25162 -1086 25210 -1058
rect 25238 -1086 25286 -1058
rect 25314 -1086 25362 -1058
rect 25390 -1086 25438 -1058
rect 25466 -1086 25522 -1058
rect 25058 -1134 25078 -1106
rect 25086 -1134 25114 -1114
rect 25162 -1134 25190 -1114
rect 25238 -1134 25266 -1114
rect 25314 -1134 25342 -1114
rect 25390 -1134 25418 -1114
rect 25466 -1134 25494 -1114
rect 25502 -1134 25522 -1106
rect 25086 -1162 25134 -1134
rect 25162 -1162 25210 -1134
rect 25238 -1162 25286 -1134
rect 25314 -1162 25362 -1134
rect 25390 -1162 25438 -1134
rect 25466 -1162 25522 -1134
rect 25058 -1210 25078 -1182
rect 25086 -1210 25114 -1190
rect 25162 -1210 25190 -1190
rect 25238 -1210 25266 -1190
rect 25314 -1210 25342 -1190
rect 25390 -1210 25418 -1190
rect 25466 -1210 25494 -1190
rect 25502 -1210 25522 -1182
rect 25086 -1238 25134 -1210
rect 25162 -1238 25210 -1210
rect 25238 -1238 25286 -1210
rect 25314 -1238 25362 -1210
rect 25390 -1238 25438 -1210
rect 25466 -1238 25522 -1210
rect 25058 -1286 25078 -1258
rect 25086 -1286 25114 -1266
rect 25162 -1286 25190 -1266
rect 25238 -1286 25266 -1266
rect 25314 -1286 25342 -1266
rect 25390 -1286 25418 -1266
rect 25466 -1286 25494 -1266
rect 25502 -1286 25522 -1258
rect 25086 -1314 25134 -1286
rect 25162 -1314 25210 -1286
rect 25238 -1314 25286 -1286
rect 25314 -1314 25362 -1286
rect 25390 -1314 25438 -1286
rect 25466 -1314 25522 -1286
rect 25058 -6118 25522 -6098
rect 25058 -6126 25078 -6118
rect 25086 -6126 25114 -6118
rect 25162 -6126 25190 -6118
rect 25238 -6126 25266 -6118
rect 25314 -6126 25342 -6118
rect 25390 -6126 25418 -6118
rect 25466 -6126 25494 -6118
rect 25502 -6126 25522 -6118
rect 25086 -6154 25134 -6126
rect 25162 -6154 25210 -6126
rect 25238 -6154 25286 -6126
rect 25314 -6154 25362 -6126
rect 25390 -6154 25438 -6126
rect 25466 -6154 25522 -6126
rect 25058 -6202 25078 -6174
rect 25086 -6202 25114 -6182
rect 25162 -6202 25190 -6182
rect 25238 -6202 25266 -6182
rect 25314 -6202 25342 -6182
rect 25390 -6202 25418 -6182
rect 25466 -6202 25494 -6182
rect 25502 -6202 25522 -6174
rect 25086 -6230 25134 -6202
rect 25162 -6230 25210 -6202
rect 25238 -6230 25286 -6202
rect 25314 -6230 25362 -6202
rect 25390 -6230 25438 -6202
rect 25466 -6230 25522 -6202
rect 25058 -6278 25078 -6250
rect 25086 -6278 25114 -6258
rect 25162 -6278 25190 -6258
rect 25238 -6278 25266 -6258
rect 25314 -6278 25342 -6258
rect 25390 -6278 25418 -6258
rect 25466 -6278 25494 -6258
rect 25502 -6278 25522 -6250
rect 25086 -6306 25134 -6278
rect 25162 -6306 25210 -6278
rect 25238 -6306 25286 -6278
rect 25314 -6306 25362 -6278
rect 25390 -6306 25438 -6278
rect 25466 -6306 25522 -6278
rect 25058 -6354 25078 -6326
rect 25086 -6354 25114 -6334
rect 25162 -6354 25190 -6334
rect 25238 -6354 25266 -6334
rect 25314 -6354 25342 -6334
rect 25390 -6354 25418 -6334
rect 25466 -6354 25494 -6334
rect 25502 -6354 25522 -6326
rect 25086 -6382 25134 -6354
rect 25162 -6382 25210 -6354
rect 25238 -6382 25286 -6354
rect 25314 -6382 25362 -6354
rect 25390 -6382 25438 -6354
rect 25466 -6382 25522 -6354
rect 25058 -6430 25078 -6402
rect 25086 -6430 25114 -6410
rect 25162 -6430 25190 -6410
rect 25238 -6430 25266 -6410
rect 25314 -6430 25342 -6410
rect 25390 -6430 25418 -6410
rect 25466 -6430 25494 -6410
rect 25502 -6430 25522 -6402
rect 25086 -6458 25134 -6430
rect 25162 -6458 25210 -6430
rect 25238 -6458 25286 -6430
rect 25314 -6458 25362 -6430
rect 25390 -6458 25438 -6430
rect 25466 -6458 25522 -6430
rect 25058 -6506 25078 -6478
rect 25086 -6506 25114 -6486
rect 25162 -6506 25190 -6486
rect 25238 -6506 25266 -6486
rect 25314 -6506 25342 -6486
rect 25390 -6506 25418 -6486
rect 25466 -6506 25494 -6486
rect 25502 -6506 25522 -6478
rect 25086 -6534 25134 -6506
rect 25162 -6534 25210 -6506
rect 25238 -6534 25286 -6506
rect 25314 -6534 25362 -6506
rect 25390 -6534 25438 -6506
rect 25466 -6534 25522 -6506
rect 24818 -7438 25282 -7418
rect 24818 -7446 24838 -7438
rect 24846 -7446 24874 -7438
rect 24922 -7446 24950 -7438
rect 24998 -7446 25026 -7438
rect 25074 -7446 25102 -7438
rect 25150 -7446 25178 -7438
rect 25226 -7446 25254 -7438
rect 25262 -7446 25282 -7438
rect 24846 -7474 24894 -7446
rect 24922 -7474 24970 -7446
rect 24998 -7474 25046 -7446
rect 25074 -7474 25122 -7446
rect 25150 -7474 25198 -7446
rect 25226 -7474 25282 -7446
rect 24818 -7522 24838 -7494
rect 24846 -7522 24874 -7502
rect 24922 -7522 24950 -7502
rect 24998 -7522 25026 -7502
rect 25074 -7522 25102 -7502
rect 25150 -7522 25178 -7502
rect 25226 -7522 25254 -7502
rect 25262 -7522 25282 -7494
rect 24846 -7550 24894 -7522
rect 24922 -7550 24970 -7522
rect 24998 -7550 25046 -7522
rect 25074 -7550 25122 -7522
rect 25150 -7550 25198 -7522
rect 25226 -7550 25282 -7522
rect 24818 -7598 24838 -7570
rect 24846 -7598 24874 -7578
rect 24922 -7598 24950 -7578
rect 24998 -7598 25026 -7578
rect 25074 -7598 25102 -7578
rect 25150 -7598 25178 -7578
rect 25226 -7598 25254 -7578
rect 25262 -7598 25282 -7570
rect 24846 -7626 24894 -7598
rect 24922 -7626 24970 -7598
rect 24998 -7626 25046 -7598
rect 25074 -7626 25122 -7598
rect 25150 -7626 25198 -7598
rect 25226 -7626 25282 -7598
rect 24818 -7674 24838 -7646
rect 24846 -7674 24874 -7654
rect 24922 -7674 24950 -7654
rect 24998 -7674 25026 -7654
rect 25074 -7674 25102 -7654
rect 25150 -7674 25178 -7654
rect 25226 -7674 25254 -7654
rect 25262 -7674 25282 -7646
rect 24846 -7702 24894 -7674
rect 24922 -7702 24970 -7674
rect 24998 -7702 25046 -7674
rect 25074 -7702 25122 -7674
rect 25150 -7702 25198 -7674
rect 25226 -7702 25282 -7674
rect 24818 -7750 24838 -7722
rect 24846 -7750 24874 -7730
rect 24922 -7750 24950 -7730
rect 24998 -7750 25026 -7730
rect 25074 -7750 25102 -7730
rect 25150 -7750 25178 -7730
rect 25226 -7750 25254 -7730
rect 25262 -7750 25282 -7722
rect 24846 -7778 24894 -7750
rect 24922 -7778 24970 -7750
rect 24998 -7778 25046 -7750
rect 25074 -7778 25122 -7750
rect 25150 -7778 25198 -7750
rect 25226 -7778 25282 -7750
rect 24818 -7826 24838 -7798
rect 24846 -7826 24874 -7806
rect 24922 -7826 24950 -7806
rect 24998 -7826 25026 -7806
rect 25074 -7826 25102 -7806
rect 25150 -7826 25178 -7806
rect 25226 -7826 25254 -7806
rect 25262 -7826 25282 -7798
rect 24846 -7840 24894 -7826
rect 24922 -7840 24970 -7826
rect 24998 -7840 25046 -7826
rect 25074 -7840 25122 -7826
rect 25150 -7840 25198 -7826
rect 25226 -7840 25282 -7826
use barth  barth_0
timestamp 1665184495
transform 1 0 5220 0 1 -3120
box -5220 -840 2940 2880
use barthmanf  barthmanf_0
timestamp 1665184495
transform 1 0 15540 0 1 -3480
box -4680 -900 7080 3060
use barthnauta  barthnauta_0
timestamp 1665184495
transform 1 0 16140 0 1 720
box -5220 -840 5340 2880
use manf  manf_0
timestamp 1665184495
transform 1 0 4680 0 1 -7200
box -4680 -900 4680 3060
use manfvieru  manfvieru_0
timestamp 1665184495
transform 1 0 29880 0 1 -11640
box -5580 -1980 16140 4500
use nauta  nauta_0
timestamp 1665184495
transform 1 0 5220 0 1 840
box -5220 -840 540 2640
use nautanauta  nautanauta_0
timestamp 1665184495
transform 1 0 29880 0 1 1860
box -5580 -1980 14940 4080
use nautavieru  nautavieru_0
timestamp 1665184495
transform 1 0 30120 0 1 -4860
box -5580 -1980 14940 4260
<< end >>
