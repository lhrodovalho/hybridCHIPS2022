magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7380 5700 -6600 6900
rect -7380 4140 -6600 5460
<< nmos >>
rect -6960 -1080 -6840 -720
<< pmos >>
rect -6960 4680 -6840 4980
<< mvpmos >>
rect -6960 6240 -6840 6600
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
<< pdiff >>
rect -7080 4883 -6960 4980
rect -7080 4837 -7043 4883
rect -6997 4837 -6960 4883
rect -7080 4763 -6960 4837
rect -7080 4717 -7043 4763
rect -6997 4717 -6960 4763
rect -7080 4680 -6960 4717
rect -6840 4883 -6720 4980
rect -6840 4837 -6803 4883
rect -6757 4837 -6720 4883
rect -6840 4763 -6720 4837
rect -6840 4717 -6803 4763
rect -6757 4717 -6720 4763
rect -6840 4680 -6720 4717
<< mvpdiff >>
rect -7080 6563 -6960 6600
rect -7080 6517 -7043 6563
rect -6997 6517 -6960 6563
rect -7080 6443 -6960 6517
rect -7080 6397 -7043 6443
rect -6997 6397 -6960 6443
rect -7080 6323 -6960 6397
rect -7080 6277 -7043 6323
rect -6997 6277 -6960 6323
rect -7080 6240 -6960 6277
rect -6840 6563 -6720 6600
rect -6840 6517 -6803 6563
rect -6757 6517 -6720 6563
rect -6840 6443 -6720 6517
rect -6840 6397 -6803 6443
rect -6757 6397 -6720 6443
rect -6840 6323 -6720 6397
rect -6840 6277 -6803 6323
rect -6757 6277 -6720 6323
rect -6840 6240 -6720 6277
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
<< pdiffc >>
rect -7043 4837 -6997 4883
rect -7043 4717 -6997 4763
rect -6803 4837 -6757 4883
rect -6803 4717 -6757 4763
<< mvpdiffc >>
rect -7043 6517 -6997 6563
rect -7043 6397 -6997 6443
rect -7043 6277 -6997 6323
rect -6803 6517 -6757 6563
rect -6803 6397 -6757 6443
rect -6803 6277 -6757 6323
<< psubdiff >>
rect -7560 7043 -6600 7080
rect -7560 6997 -7523 7043
rect -7477 6997 -7403 7043
rect -7357 6997 -7283 7043
rect -7237 6997 -7163 7043
rect -7117 6997 -7043 7043
rect -6997 6997 -6923 7043
rect -6877 6997 -6803 7043
rect -6757 6997 -6683 7043
rect -6637 6997 -6600 7043
rect -7560 6960 -6600 6997
rect -7560 6923 -7440 6960
rect -7560 6877 -7523 6923
rect -7477 6877 -7440 6923
rect -7560 6803 -7440 6877
rect -7560 6757 -7523 6803
rect -7477 6757 -7440 6803
rect -7560 6683 -7440 6757
rect -7560 6637 -7523 6683
rect -7477 6637 -7440 6683
rect -7560 6563 -7440 6637
rect -7560 6517 -7523 6563
rect -7477 6517 -7440 6563
rect -7560 6443 -7440 6517
rect -7560 6397 -7523 6443
rect -7477 6397 -7440 6443
rect -7560 6323 -7440 6397
rect -7560 6277 -7523 6323
rect -7477 6277 -7440 6323
rect -7560 6203 -7440 6277
rect -7560 6157 -7523 6203
rect -7477 6157 -7440 6203
rect -7560 6083 -7440 6157
rect -7560 6037 -7523 6083
rect -7477 6037 -7440 6083
rect -7560 5963 -7440 6037
rect -7560 5917 -7523 5963
rect -7477 5917 -7440 5963
rect -7560 5843 -7440 5917
rect -7560 5797 -7523 5843
rect -7477 5797 -7440 5843
rect -7560 5723 -7440 5797
rect -7560 5677 -7523 5723
rect -7477 5677 -7440 5723
rect -7560 5640 -7440 5677
rect -7560 5603 -6600 5640
rect -7560 5557 -7523 5603
rect -7477 5557 -7403 5603
rect -7357 5557 -7283 5603
rect -7237 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6600 5603
rect -7560 5520 -6600 5557
rect -7560 5483 -7440 5520
rect -7560 5437 -7523 5483
rect -7477 5437 -7440 5483
rect -7560 5363 -7440 5437
rect -7560 5317 -7523 5363
rect -7477 5317 -7440 5363
rect -7560 5243 -7440 5317
rect -7560 5197 -7523 5243
rect -7477 5197 -7440 5243
rect -7560 5123 -7440 5197
rect -7560 5077 -7523 5123
rect -7477 5077 -7440 5123
rect -7560 5003 -7440 5077
rect -7560 4957 -7523 5003
rect -7477 4957 -7440 5003
rect -7560 4883 -7440 4957
rect -7560 4837 -7523 4883
rect -7477 4837 -7440 4883
rect -7560 4763 -7440 4837
rect -7560 4717 -7523 4763
rect -7477 4717 -7440 4763
rect -7560 4643 -7440 4717
rect -7560 4597 -7523 4643
rect -7477 4597 -7440 4643
rect -7560 4523 -7440 4597
rect -7560 4477 -7523 4523
rect -7477 4477 -7440 4523
rect -7560 4403 -7440 4477
rect -7560 4357 -7523 4403
rect -7477 4357 -7440 4403
rect -7560 4283 -7440 4357
rect -7560 4237 -7523 4283
rect -7477 4237 -7440 4283
rect -7560 4163 -7440 4237
rect -7560 4117 -7523 4163
rect -7477 4117 -7440 4163
rect -7560 4080 -7440 4117
rect -7560 4043 -6600 4080
rect -7560 3997 -7523 4043
rect -7477 3997 -7403 4043
rect -7357 3997 -7283 4043
rect -7237 3997 -7163 4043
rect -7117 3997 -7043 4043
rect -6997 3997 -6923 4043
rect -6877 3997 -6803 4043
rect -6757 3997 -6683 4043
rect -6637 3997 -6600 4043
rect -7560 3960 -6600 3997
rect -7560 3923 -7440 3960
rect -7560 3877 -7523 3923
rect -7477 3877 -7440 3923
rect -7560 3803 -7440 3877
rect -7560 3757 -7523 3803
rect -7477 3757 -7440 3803
rect -7560 3563 -7440 3757
rect -7560 3517 -7523 3563
rect -7477 3517 -7440 3563
rect -7560 3443 -7440 3517
rect -7560 3397 -7523 3443
rect -7477 3397 -7440 3443
rect -7560 3323 -7440 3397
rect -7560 3277 -7523 3323
rect -7477 3277 -7440 3323
rect -7560 3083 -7440 3277
rect -7560 3037 -7523 3083
rect -7477 3037 -7440 3083
rect -7560 2963 -7440 3037
rect -7560 2917 -7523 2963
rect -7477 2917 -7440 2963
rect -7560 2880 -7440 2917
rect -7560 2843 -6600 2880
rect -7560 2797 -7523 2843
rect -7477 2797 -7403 2843
rect -7357 2797 -7283 2843
rect -7237 2797 -7163 2843
rect -7117 2797 -7043 2843
rect -6997 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6683 2843
rect -6637 2797 -6600 2843
rect -7560 2760 -6600 2797
rect -7560 2723 -7440 2760
rect -7560 2677 -7523 2723
rect -7477 2677 -7440 2723
rect -7560 2603 -7440 2677
rect -7560 2557 -7523 2603
rect -7477 2557 -7440 2603
rect -7560 2483 -7440 2557
rect -7560 2437 -7523 2483
rect -7477 2437 -7440 2483
rect -7560 2400 -7440 2437
rect -7560 2363 -6600 2400
rect -7560 2317 -7523 2363
rect -7477 2317 -7403 2363
rect -7357 2317 -7283 2363
rect -7237 2317 -7163 2363
rect -7117 2317 -7043 2363
rect -6997 2317 -6923 2363
rect -6877 2317 -6803 2363
rect -6757 2317 -6683 2363
rect -6637 2317 -6600 2363
rect -7560 2280 -6600 2317
rect -7560 2243 -7440 2280
rect -7560 2197 -7523 2243
rect -7477 2197 -7440 2243
rect -7560 2123 -7440 2197
rect -7560 2077 -7523 2123
rect -7477 2077 -7440 2123
rect -7560 2003 -7440 2077
rect -7560 1957 -7523 2003
rect -7477 1957 -7440 2003
rect -7560 1920 -7440 1957
rect -7560 1883 -6600 1920
rect -7560 1837 -7523 1883
rect -7477 1837 -7403 1883
rect -7357 1837 -7283 1883
rect -7237 1837 -7163 1883
rect -7117 1837 -7043 1883
rect -6997 1837 -6923 1883
rect -6877 1837 -6803 1883
rect -6757 1837 -6683 1883
rect -6637 1837 -6600 1883
rect -7560 1800 -6600 1837
rect -7560 1763 -7440 1800
rect -7560 1717 -7523 1763
rect -7477 1717 -7440 1763
rect -7560 1643 -7440 1717
rect -7560 1597 -7523 1643
rect -7477 1597 -7440 1643
rect -7560 1523 -7440 1597
rect -7560 1477 -7523 1523
rect -7477 1477 -7440 1523
rect -7560 1440 -7440 1477
rect -7560 1403 -6600 1440
rect -7560 1357 -7523 1403
rect -7477 1357 -7403 1403
rect -7357 1357 -7283 1403
rect -7237 1357 -7163 1403
rect -7117 1357 -7043 1403
rect -6997 1357 -6923 1403
rect -6877 1357 -6803 1403
rect -6757 1357 -6683 1403
rect -6637 1357 -6600 1403
rect -7560 1320 -6600 1357
rect -7560 1283 -7440 1320
rect -7560 1237 -7523 1283
rect -7477 1237 -7440 1283
rect -7560 1163 -7440 1237
rect -7560 1117 -7523 1163
rect -7477 1117 -7440 1163
rect -7560 1043 -7440 1117
rect -7560 997 -7523 1043
rect -7477 997 -7440 1043
rect -7560 960 -7440 997
rect -7560 923 -6600 960
rect -7560 877 -7523 923
rect -7477 877 -7403 923
rect -7357 877 -7283 923
rect -7237 877 -7163 923
rect -7117 877 -7043 923
rect -6997 877 -6923 923
rect -6877 877 -6803 923
rect -6757 877 -6683 923
rect -6637 877 -6600 923
rect -7560 840 -6600 877
rect -7560 803 -7440 840
rect -7560 757 -7523 803
rect -7477 757 -7440 803
rect -7560 683 -7440 757
rect -7560 637 -7523 683
rect -7477 637 -7440 683
rect -7560 443 -7440 637
rect -7560 397 -7523 443
rect -7477 397 -7440 443
rect -7560 323 -7440 397
rect -7560 277 -7523 323
rect -7477 277 -7440 323
rect -7560 203 -7440 277
rect -7560 157 -7523 203
rect -7477 157 -7440 203
rect -7560 -37 -7440 157
rect -7560 -83 -7523 -37
rect -7477 -83 -7440 -37
rect -7560 -157 -7440 -83
rect -7560 -203 -7523 -157
rect -7477 -203 -7440 -157
rect -7560 -240 -7440 -203
rect -7560 -277 -6600 -240
rect -7560 -323 -7523 -277
rect -7477 -323 -7403 -277
rect -7357 -323 -7283 -277
rect -7237 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6600 -277
rect -7560 -360 -6600 -323
rect -7560 -397 -7440 -360
rect -7560 -443 -7523 -397
rect -7477 -443 -7440 -397
rect -7560 -517 -7440 -443
rect -7560 -563 -7523 -517
rect -7477 -563 -7440 -517
rect -7560 -637 -7440 -563
rect -7560 -683 -7523 -637
rect -7477 -683 -7440 -637
rect -7560 -757 -7440 -683
rect -7560 -803 -7523 -757
rect -7477 -803 -7440 -757
rect -7560 -877 -7440 -803
rect -7560 -923 -7523 -877
rect -7477 -923 -7440 -877
rect -7560 -997 -7440 -923
rect -7560 -1043 -7523 -997
rect -7477 -1043 -7440 -997
rect -7560 -1117 -7440 -1043
rect -7560 -1163 -7523 -1117
rect -7477 -1163 -7440 -1117
rect -7560 -1200 -7440 -1163
rect -7560 -1237 -6600 -1200
rect -7560 -1283 -7523 -1237
rect -7477 -1283 -7403 -1237
rect -7357 -1283 -7283 -1237
rect -7237 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6600 -1237
rect -7560 -1320 -6600 -1283
<< nsubdiff >>
rect -7320 5363 -6720 5400
rect -7320 5317 -7283 5363
rect -7237 5317 -7163 5363
rect -7117 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6720 5363
rect -7320 5280 -6720 5317
rect -7320 5243 -7200 5280
rect -7320 5197 -7283 5243
rect -7237 5197 -7200 5243
rect -7320 5123 -7200 5197
rect -7320 5077 -7283 5123
rect -7237 5077 -7200 5123
rect -7320 5003 -7200 5077
rect -7320 4957 -7283 5003
rect -7237 4957 -7200 5003
rect -7320 4883 -7200 4957
rect -7320 4837 -7283 4883
rect -7237 4837 -7200 4883
rect -7320 4763 -7200 4837
rect -7320 4717 -7283 4763
rect -7237 4717 -7200 4763
rect -7320 4643 -7200 4717
rect -7320 4597 -7283 4643
rect -7237 4597 -7200 4643
rect -7320 4523 -7200 4597
rect -7320 4477 -7283 4523
rect -7237 4477 -7200 4523
rect -7320 4403 -7200 4477
rect -7320 4357 -7283 4403
rect -7237 4357 -7200 4403
rect -7320 4320 -7200 4357
rect -7320 4283 -6720 4320
rect -7320 4237 -7283 4283
rect -7237 4237 -7163 4283
rect -7117 4237 -7043 4283
rect -6997 4237 -6923 4283
rect -6877 4237 -6803 4283
rect -6757 4237 -6720 4283
rect -7320 4200 -6720 4237
<< mvnsubdiff >>
rect -7320 6803 -6720 6840
rect -7320 6757 -7283 6803
rect -7237 6757 -7163 6803
rect -7117 6757 -7043 6803
rect -6997 6757 -6923 6803
rect -6877 6757 -6803 6803
rect -6757 6757 -6720 6803
rect -7320 6720 -6720 6757
rect -7320 6683 -7200 6720
rect -7320 6637 -7283 6683
rect -7237 6637 -7200 6683
rect -7320 6563 -7200 6637
rect -7320 6517 -7283 6563
rect -7237 6517 -7200 6563
rect -7320 6443 -7200 6517
rect -7320 6397 -7283 6443
rect -7237 6397 -7200 6443
rect -7320 6323 -7200 6397
rect -7320 6277 -7283 6323
rect -7237 6277 -7200 6323
rect -7320 6203 -7200 6277
rect -7320 6157 -7283 6203
rect -7237 6157 -7200 6203
rect -7320 6083 -7200 6157
rect -7320 6037 -7283 6083
rect -7237 6037 -7200 6083
rect -7320 5963 -7200 6037
rect -7320 5917 -7283 5963
rect -7237 5917 -7200 5963
rect -7320 5880 -7200 5917
rect -7320 5843 -6720 5880
rect -7320 5797 -7283 5843
rect -7237 5797 -7163 5843
rect -7117 5797 -7043 5843
rect -6997 5797 -6923 5843
rect -6877 5797 -6803 5843
rect -6757 5797 -6720 5843
rect -7320 5760 -6720 5797
<< psubdiffcont >>
rect -7523 6997 -7477 7043
rect -7403 6997 -7357 7043
rect -7283 6997 -7237 7043
rect -7163 6997 -7117 7043
rect -7043 6997 -6997 7043
rect -6923 6997 -6877 7043
rect -6803 6997 -6757 7043
rect -6683 6997 -6637 7043
rect -7523 6877 -7477 6923
rect -7523 6757 -7477 6803
rect -7523 6637 -7477 6683
rect -7523 6517 -7477 6563
rect -7523 6397 -7477 6443
rect -7523 6277 -7477 6323
rect -7523 6157 -7477 6203
rect -7523 6037 -7477 6083
rect -7523 5917 -7477 5963
rect -7523 5797 -7477 5843
rect -7523 5677 -7477 5723
rect -7523 5557 -7477 5603
rect -7403 5557 -7357 5603
rect -7283 5557 -7237 5603
rect -7163 5557 -7117 5603
rect -7043 5557 -6997 5603
rect -6923 5557 -6877 5603
rect -6803 5557 -6757 5603
rect -6683 5557 -6637 5603
rect -7523 5437 -7477 5483
rect -7523 5317 -7477 5363
rect -7523 5197 -7477 5243
rect -7523 5077 -7477 5123
rect -7523 4957 -7477 5003
rect -7523 4837 -7477 4883
rect -7523 4717 -7477 4763
rect -7523 4597 -7477 4643
rect -7523 4477 -7477 4523
rect -7523 4357 -7477 4403
rect -7523 4237 -7477 4283
rect -7523 4117 -7477 4163
rect -7523 3997 -7477 4043
rect -7403 3997 -7357 4043
rect -7283 3997 -7237 4043
rect -7163 3997 -7117 4043
rect -7043 3997 -6997 4043
rect -6923 3997 -6877 4043
rect -6803 3997 -6757 4043
rect -6683 3997 -6637 4043
rect -7523 3877 -7477 3923
rect -7523 3757 -7477 3803
rect -7523 3517 -7477 3563
rect -7523 3397 -7477 3443
rect -7523 3277 -7477 3323
rect -7523 3037 -7477 3083
rect -7523 2917 -7477 2963
rect -7523 2797 -7477 2843
rect -7403 2797 -7357 2843
rect -7283 2797 -7237 2843
rect -7163 2797 -7117 2843
rect -7043 2797 -6997 2843
rect -6923 2797 -6877 2843
rect -6803 2797 -6757 2843
rect -6683 2797 -6637 2843
rect -7523 2677 -7477 2723
rect -7523 2557 -7477 2603
rect -7523 2437 -7477 2483
rect -7523 2317 -7477 2363
rect -7403 2317 -7357 2363
rect -7283 2317 -7237 2363
rect -7163 2317 -7117 2363
rect -7043 2317 -6997 2363
rect -6923 2317 -6877 2363
rect -6803 2317 -6757 2363
rect -6683 2317 -6637 2363
rect -7523 2197 -7477 2243
rect -7523 2077 -7477 2123
rect -7523 1957 -7477 2003
rect -7523 1837 -7477 1883
rect -7403 1837 -7357 1883
rect -7283 1837 -7237 1883
rect -7163 1837 -7117 1883
rect -7043 1837 -6997 1883
rect -6923 1837 -6877 1883
rect -6803 1837 -6757 1883
rect -6683 1837 -6637 1883
rect -7523 1717 -7477 1763
rect -7523 1597 -7477 1643
rect -7523 1477 -7477 1523
rect -7523 1357 -7477 1403
rect -7403 1357 -7357 1403
rect -7283 1357 -7237 1403
rect -7163 1357 -7117 1403
rect -7043 1357 -6997 1403
rect -6923 1357 -6877 1403
rect -6803 1357 -6757 1403
rect -6683 1357 -6637 1403
rect -7523 1237 -7477 1283
rect -7523 1117 -7477 1163
rect -7523 997 -7477 1043
rect -7523 877 -7477 923
rect -7403 877 -7357 923
rect -7283 877 -7237 923
rect -7163 877 -7117 923
rect -7043 877 -6997 923
rect -6923 877 -6877 923
rect -6803 877 -6757 923
rect -6683 877 -6637 923
rect -7523 757 -7477 803
rect -7523 637 -7477 683
rect -7523 397 -7477 443
rect -7523 277 -7477 323
rect -7523 157 -7477 203
rect -7523 -83 -7477 -37
rect -7523 -203 -7477 -157
rect -7523 -323 -7477 -277
rect -7403 -323 -7357 -277
rect -7283 -323 -7237 -277
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -7523 -443 -7477 -397
rect -7523 -563 -7477 -517
rect -7523 -683 -7477 -637
rect -7523 -803 -7477 -757
rect -7523 -923 -7477 -877
rect -7523 -1043 -7477 -997
rect -7523 -1163 -7477 -1117
rect -7523 -1283 -7477 -1237
rect -7403 -1283 -7357 -1237
rect -7283 -1283 -7237 -1237
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
<< nsubdiffcont >>
rect -7283 5317 -7237 5363
rect -7163 5317 -7117 5363
rect -7043 5317 -6997 5363
rect -6923 5317 -6877 5363
rect -6803 5317 -6757 5363
rect -7283 5197 -7237 5243
rect -7283 5077 -7237 5123
rect -7283 4957 -7237 5003
rect -7283 4837 -7237 4883
rect -7283 4717 -7237 4763
rect -7283 4597 -7237 4643
rect -7283 4477 -7237 4523
rect -7283 4357 -7237 4403
rect -7283 4237 -7237 4283
rect -7163 4237 -7117 4283
rect -7043 4237 -6997 4283
rect -6923 4237 -6877 4283
rect -6803 4237 -6757 4283
<< mvnsubdiffcont >>
rect -7283 6757 -7237 6803
rect -7163 6757 -7117 6803
rect -7043 6757 -6997 6803
rect -6923 6757 -6877 6803
rect -6803 6757 -6757 6803
rect -7283 6637 -7237 6683
rect -7283 6517 -7237 6563
rect -7283 6397 -7237 6443
rect -7283 6277 -7237 6323
rect -7283 6157 -7237 6203
rect -7283 6037 -7237 6083
rect -7283 5917 -7237 5963
rect -7283 5797 -7237 5843
rect -7163 5797 -7117 5843
rect -7043 5797 -6997 5843
rect -6923 5797 -6877 5843
rect -6803 5797 -6757 5843
<< polysilicon >>
rect -6960 6600 -6840 6660
rect -6960 6083 -6840 6240
rect -6960 6037 -6923 6083
rect -6877 6037 -6840 6083
rect -6960 6000 -6840 6037
rect -6960 4980 -6840 5040
rect -6960 4523 -6840 4680
rect -6960 4477 -6923 4523
rect -6877 4477 -6840 4523
rect -6960 4440 -6840 4477
rect -6960 -517 -6840 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6840 -517
rect -6960 -720 -6840 -563
rect -6960 -1140 -6840 -1080
<< polycontact >>
rect -6923 6037 -6877 6083
rect -6923 4477 -6877 4523
rect -6923 -563 -6877 -517
<< metal1 >>
rect -7560 7043 -6600 7080
rect -7560 6997 -7523 7043
rect -7477 6997 -7403 7043
rect -7357 6997 -7283 7043
rect -7237 6997 -7163 7043
rect -7117 6997 -7043 7043
rect -6997 6997 -6923 7043
rect -6877 6997 -6803 7043
rect -6757 6997 -6683 7043
rect -6637 6997 -6600 7043
rect -7560 6960 -6600 6997
rect -7560 6923 -7440 6960
rect -7560 6877 -7523 6923
rect -7477 6877 -7440 6923
rect -7560 6803 -7440 6877
rect -7560 6757 -7523 6803
rect -7477 6757 -7440 6803
rect -7560 6683 -7440 6757
rect -7560 6637 -7523 6683
rect -7477 6637 -7440 6683
rect -7560 6563 -7440 6637
rect -7560 6517 -7523 6563
rect -7477 6517 -7440 6563
rect -7560 6443 -7440 6517
rect -7560 6397 -7523 6443
rect -7477 6397 -7440 6443
rect -7560 6323 -7440 6397
rect -7560 6277 -7523 6323
rect -7477 6277 -7440 6323
rect -7560 6203 -7440 6277
rect -7560 6157 -7523 6203
rect -7477 6157 -7440 6203
rect -7560 6083 -7440 6157
rect -7560 6037 -7523 6083
rect -7477 6037 -7440 6083
rect -7560 5963 -7440 6037
rect -7560 5917 -7523 5963
rect -7477 5917 -7440 5963
rect -7560 5843 -7440 5917
rect -7560 5797 -7523 5843
rect -7477 5797 -7440 5843
rect -7560 5723 -7440 5797
rect -7320 6806 -6600 6840
rect -7320 6803 -6806 6806
rect -7320 6757 -7283 6803
rect -7237 6757 -7163 6803
rect -7117 6757 -7043 6803
rect -6997 6757 -6923 6803
rect -6877 6757 -6806 6803
rect -7320 6754 -6806 6757
rect -6754 6754 -6600 6806
rect -7320 6720 -6600 6754
rect -7320 6683 -7200 6720
rect -7320 6637 -7283 6683
rect -7237 6637 -7200 6683
rect -7320 6563 -7200 6637
rect -7320 6517 -7283 6563
rect -7237 6517 -7200 6563
rect -7320 6443 -7200 6517
rect -7320 6397 -7283 6443
rect -7237 6397 -7200 6443
rect -7320 6323 -7200 6397
rect -7320 6277 -7283 6323
rect -7237 6277 -7200 6323
rect -7320 6203 -7200 6277
rect -7320 6157 -7283 6203
rect -7237 6157 -7200 6203
rect -7320 6083 -7200 6157
rect -7320 6037 -7283 6083
rect -7237 6037 -7200 6083
rect -7320 5963 -7200 6037
rect -7080 6563 -6960 6600
rect -7080 6517 -7043 6563
rect -6997 6517 -6960 6563
rect -7080 6443 -6960 6517
rect -7080 6397 -7043 6443
rect -6997 6397 -6960 6443
rect -7080 6323 -6960 6397
rect -7080 6277 -7043 6323
rect -6997 6277 -6960 6323
rect -7080 6120 -6960 6277
rect -6840 6566 -6720 6600
rect -6840 6514 -6806 6566
rect -6754 6514 -6720 6566
rect -6840 6446 -6720 6514
rect -6840 6394 -6806 6446
rect -6754 6394 -6720 6446
rect -6840 6326 -6720 6394
rect -6840 6274 -6806 6326
rect -6754 6274 -6720 6326
rect -6840 6240 -6720 6274
rect -7080 6083 -6840 6120
rect -7080 6037 -6923 6083
rect -6877 6037 -6840 6083
rect -7080 6000 -6840 6037
rect -7320 5917 -7283 5963
rect -7237 5917 -7200 5963
rect -7320 5880 -7200 5917
rect -7320 5843 -6600 5880
rect -7320 5797 -7283 5843
rect -7237 5797 -7163 5843
rect -7117 5797 -7043 5843
rect -6997 5797 -6923 5843
rect -6877 5797 -6803 5843
rect -6757 5797 -6600 5843
rect -7320 5760 -6600 5797
rect -7560 5677 -7523 5723
rect -7477 5677 -7440 5723
rect -7560 5640 -7440 5677
rect -7560 5603 -6600 5640
rect -7560 5557 -7523 5603
rect -7477 5557 -7403 5603
rect -7357 5557 -7283 5603
rect -7237 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6600 5603
rect -7560 5520 -6600 5557
rect -7560 5483 -7440 5520
rect -7560 5437 -7523 5483
rect -7477 5437 -7440 5483
rect -7560 5363 -7440 5437
rect -7560 5317 -7523 5363
rect -7477 5317 -7440 5363
rect -7560 5243 -7440 5317
rect -7560 5197 -7523 5243
rect -7477 5197 -7440 5243
rect -7560 5123 -7440 5197
rect -7560 5077 -7523 5123
rect -7477 5077 -7440 5123
rect -7560 5003 -7440 5077
rect -7560 4957 -7523 5003
rect -7477 4957 -7440 5003
rect -7560 4883 -7440 4957
rect -7560 4837 -7523 4883
rect -7477 4837 -7440 4883
rect -7560 4763 -7440 4837
rect -7560 4717 -7523 4763
rect -7477 4717 -7440 4763
rect -7560 4643 -7440 4717
rect -7560 4597 -7523 4643
rect -7477 4597 -7440 4643
rect -7560 4523 -7440 4597
rect -7560 4477 -7523 4523
rect -7477 4477 -7440 4523
rect -7560 4403 -7440 4477
rect -7560 4357 -7523 4403
rect -7477 4357 -7440 4403
rect -7560 4283 -7440 4357
rect -7560 4237 -7523 4283
rect -7477 4237 -7440 4283
rect -7560 4163 -7440 4237
rect -7320 5363 -6720 5400
rect -7320 5317 -7283 5363
rect -7237 5317 -7163 5363
rect -7117 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6720 5363
rect -7320 5280 -6720 5317
rect -7320 5243 -7200 5280
rect -7320 5197 -7283 5243
rect -7237 5197 -7200 5243
rect -7320 5123 -7200 5197
rect -7320 5077 -7283 5123
rect -7237 5077 -7200 5123
rect -7320 5003 -7200 5077
rect -7320 4957 -7283 5003
rect -7237 4957 -7200 5003
rect -7320 4883 -7200 4957
rect -7320 4837 -7283 4883
rect -7237 4837 -7200 4883
rect -7320 4763 -7200 4837
rect -7320 4717 -7283 4763
rect -7237 4717 -7200 4763
rect -7320 4643 -7200 4717
rect -7320 4597 -7283 4643
rect -7237 4597 -7200 4643
rect -7320 4523 -7200 4597
rect -7320 4477 -7283 4523
rect -7237 4477 -7200 4523
rect -7320 4403 -7200 4477
rect -7080 4883 -6960 4980
rect -7080 4837 -7043 4883
rect -6997 4837 -6960 4883
rect -7080 4763 -6960 4837
rect -7080 4717 -7043 4763
rect -6997 4717 -6960 4763
rect -7080 4560 -6960 4717
rect -6840 4886 -6720 4980
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4766 -6720 4834
rect -6840 4714 -6806 4766
rect -6754 4714 -6720 4766
rect -6840 4680 -6720 4714
rect -7080 4523 -6840 4560
rect -7080 4477 -6923 4523
rect -6877 4477 -6840 4523
rect -7080 4440 -6840 4477
rect -7320 4357 -7283 4403
rect -7237 4357 -7200 4403
rect -7320 4320 -7200 4357
rect -7320 4286 -6600 4320
rect -7320 4234 -7286 4286
rect -7234 4283 -6600 4286
rect -7234 4237 -7163 4283
rect -7117 4237 -7043 4283
rect -6997 4237 -6923 4283
rect -6877 4237 -6803 4283
rect -6757 4237 -6600 4283
rect -7234 4234 -6600 4237
rect -7320 4200 -6600 4234
rect -7560 4117 -7523 4163
rect -7477 4117 -7440 4163
rect -7560 4080 -7440 4117
rect -7560 4046 -6600 4080
rect -7560 4043 -6806 4046
rect -6754 4043 -6600 4046
rect -7560 3997 -7523 4043
rect -7477 3997 -7403 4043
rect -7357 3997 -7283 4043
rect -7237 3997 -7163 4043
rect -7117 3997 -7043 4043
rect -6997 3997 -6923 4043
rect -6877 3997 -6806 4043
rect -6754 3997 -6683 4043
rect -6637 3997 -6600 4043
rect -7560 3994 -6806 3997
rect -6754 3994 -6600 3997
rect -7560 3960 -6600 3994
rect -7560 3923 -7440 3960
rect -7560 3877 -7523 3923
rect -7477 3877 -7440 3923
rect -7560 3803 -7440 3877
rect -7560 3757 -7523 3803
rect -7477 3757 -7440 3803
rect -7560 3563 -7440 3757
rect -7560 3517 -7523 3563
rect -7477 3517 -7440 3563
rect -7560 3443 -7440 3517
rect -7560 3397 -7523 3443
rect -7477 3397 -7440 3443
rect -7560 3323 -7440 3397
rect -7560 3277 -7523 3323
rect -7477 3277 -7440 3323
rect -7560 3083 -7440 3277
rect -7560 3037 -7523 3083
rect -7477 3037 -7440 3083
rect -7560 2963 -7440 3037
rect -7560 2917 -7523 2963
rect -7477 2917 -7440 2963
rect -7560 2880 -7440 2917
rect -7560 2846 -6600 2880
rect -7560 2843 -6806 2846
rect -6754 2843 -6600 2846
rect -7560 2797 -7523 2843
rect -7477 2797 -7403 2843
rect -7357 2797 -7283 2843
rect -7237 2797 -7163 2843
rect -7117 2797 -7043 2843
rect -6997 2797 -6923 2843
rect -6877 2797 -6806 2843
rect -6754 2797 -6683 2843
rect -6637 2797 -6600 2843
rect -7560 2794 -6806 2797
rect -6754 2794 -6600 2797
rect -7560 2760 -6600 2794
rect -7560 2723 -7440 2760
rect -7560 2677 -7523 2723
rect -7477 2677 -7440 2723
rect -7560 2603 -7440 2677
rect -7560 2557 -7523 2603
rect -7477 2557 -7440 2603
rect -7560 2483 -7440 2557
rect -7560 2437 -7523 2483
rect -7477 2437 -7440 2483
rect -7560 2400 -7440 2437
rect -7560 2366 -6600 2400
rect -7560 2363 -6806 2366
rect -6754 2363 -6600 2366
rect -7560 2317 -7523 2363
rect -7477 2317 -7403 2363
rect -7357 2317 -7283 2363
rect -7237 2317 -7163 2363
rect -7117 2317 -7043 2363
rect -6997 2317 -6923 2363
rect -6877 2317 -6806 2363
rect -6754 2317 -6683 2363
rect -6637 2317 -6600 2363
rect -7560 2314 -6806 2317
rect -6754 2314 -6600 2317
rect -7560 2280 -6600 2314
rect -7560 2243 -7440 2280
rect -7560 2197 -7523 2243
rect -7477 2197 -7440 2243
rect -7560 2123 -7440 2197
rect -7560 2077 -7523 2123
rect -7477 2077 -7440 2123
rect -7560 2003 -7440 2077
rect -7560 1957 -7523 2003
rect -7477 1957 -7440 2003
rect -7560 1920 -7440 1957
rect -7560 1886 -6600 1920
rect -7560 1883 -6806 1886
rect -6754 1883 -6600 1886
rect -7560 1837 -7523 1883
rect -7477 1837 -7403 1883
rect -7357 1837 -7283 1883
rect -7237 1837 -7163 1883
rect -7117 1837 -7043 1883
rect -6997 1837 -6923 1883
rect -6877 1837 -6806 1883
rect -6754 1837 -6683 1883
rect -6637 1837 -6600 1883
rect -7560 1834 -6806 1837
rect -6754 1834 -6600 1837
rect -7560 1800 -6600 1834
rect -7560 1763 -7440 1800
rect -7560 1717 -7523 1763
rect -7477 1717 -7440 1763
rect -7560 1643 -7440 1717
rect -7560 1597 -7523 1643
rect -7477 1597 -7440 1643
rect -7560 1523 -7440 1597
rect -7560 1477 -7523 1523
rect -7477 1477 -7440 1523
rect -7560 1440 -7440 1477
rect -7560 1406 -6600 1440
rect -7560 1403 -6806 1406
rect -6754 1403 -6600 1406
rect -7560 1357 -7523 1403
rect -7477 1357 -7403 1403
rect -7357 1357 -7283 1403
rect -7237 1357 -7163 1403
rect -7117 1357 -7043 1403
rect -6997 1357 -6923 1403
rect -6877 1357 -6806 1403
rect -6754 1357 -6683 1403
rect -6637 1357 -6600 1403
rect -7560 1354 -6806 1357
rect -6754 1354 -6600 1357
rect -7560 1320 -6600 1354
rect -7560 1283 -7440 1320
rect -7560 1237 -7523 1283
rect -7477 1237 -7440 1283
rect -7560 1163 -7440 1237
rect -7560 1117 -7523 1163
rect -7477 1117 -7440 1163
rect -7560 1043 -7440 1117
rect -7560 997 -7523 1043
rect -7477 997 -7440 1043
rect -7560 960 -7440 997
rect -7560 926 -6600 960
rect -7560 923 -6806 926
rect -6754 923 -6600 926
rect -7560 877 -7523 923
rect -7477 877 -7403 923
rect -7357 877 -7283 923
rect -7237 877 -7163 923
rect -7117 877 -7043 923
rect -6997 877 -6923 923
rect -6877 877 -6806 923
rect -6754 877 -6683 923
rect -6637 877 -6600 923
rect -7560 874 -6806 877
rect -6754 874 -6600 877
rect -7560 840 -6600 874
rect -7560 803 -7440 840
rect -7560 757 -7523 803
rect -7477 757 -7440 803
rect -7560 683 -7440 757
rect -7560 637 -7523 683
rect -7477 637 -7440 683
rect -7560 443 -7440 637
rect -7560 397 -7523 443
rect -7477 397 -7440 443
rect -7560 323 -7440 397
rect -7560 277 -7523 323
rect -7477 277 -7440 323
rect -7560 203 -7440 277
rect -7560 157 -7523 203
rect -7477 157 -7440 203
rect -7560 -37 -7440 157
rect -7560 -83 -7523 -37
rect -7477 -83 -7440 -37
rect -7560 -157 -7440 -83
rect -7560 -203 -7523 -157
rect -7477 -203 -7440 -157
rect -7560 -240 -7440 -203
rect -7560 -274 -6600 -240
rect -7560 -277 -6806 -274
rect -6754 -277 -6600 -274
rect -7560 -323 -7523 -277
rect -7477 -323 -7403 -277
rect -7357 -323 -7283 -277
rect -7237 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6806 -277
rect -6754 -323 -6683 -277
rect -6637 -323 -6600 -277
rect -7560 -326 -6806 -323
rect -6754 -326 -6600 -323
rect -7560 -360 -6600 -326
rect -7560 -397 -7440 -360
rect -7560 -443 -7523 -397
rect -7477 -443 -7440 -397
rect -7560 -517 -7440 -443
rect -7560 -563 -7523 -517
rect -7477 -563 -7440 -517
rect -7560 -637 -7440 -563
rect -7560 -683 -7523 -637
rect -7477 -683 -7440 -637
rect -7560 -757 -7440 -683
rect -7560 -803 -7523 -757
rect -7477 -803 -7440 -757
rect -7560 -877 -7440 -803
rect -7560 -923 -7523 -877
rect -7477 -923 -7440 -877
rect -7560 -997 -7440 -923
rect -7560 -1043 -7523 -997
rect -7477 -1043 -7440 -997
rect -7560 -1117 -7440 -1043
rect -7080 -517 -6840 -480
rect -7080 -563 -6923 -517
rect -6877 -563 -6840 -517
rect -7080 -600 -6840 -563
rect -7080 -757 -6960 -600
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -754 -6720 -720
rect -6840 -806 -6806 -754
rect -6754 -806 -6720 -754
rect -6840 -874 -6720 -806
rect -6840 -926 -6806 -874
rect -6754 -926 -6720 -874
rect -6840 -994 -6720 -926
rect -6840 -1046 -6806 -994
rect -6754 -1046 -6720 -994
rect -6840 -1080 -6720 -1046
rect -7560 -1163 -7523 -1117
rect -7477 -1163 -7440 -1117
rect -7560 -1200 -7440 -1163
rect -7560 -1234 -6600 -1200
rect -7560 -1237 -6806 -1234
rect -6754 -1237 -6600 -1234
rect -7560 -1283 -7523 -1237
rect -7477 -1283 -7403 -1237
rect -7357 -1283 -7283 -1237
rect -7237 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6806 -1237
rect -6754 -1283 -6683 -1237
rect -6637 -1283 -6600 -1237
rect -7560 -1286 -6806 -1283
rect -6754 -1286 -6600 -1283
rect -7560 -1320 -6600 -1286
<< via1 >>
rect -6806 6803 -6754 6806
rect -6806 6757 -6803 6803
rect -6803 6757 -6757 6803
rect -6757 6757 -6754 6803
rect -6806 6754 -6754 6757
rect -6806 6563 -6754 6566
rect -6806 6517 -6803 6563
rect -6803 6517 -6757 6563
rect -6757 6517 -6754 6563
rect -6806 6514 -6754 6517
rect -6806 6443 -6754 6446
rect -6806 6397 -6803 6443
rect -6803 6397 -6757 6443
rect -6757 6397 -6754 6443
rect -6806 6394 -6754 6397
rect -6806 6323 -6754 6326
rect -6806 6277 -6803 6323
rect -6803 6277 -6757 6323
rect -6757 6277 -6754 6323
rect -6806 6274 -6754 6277
rect -6806 4883 -6754 4886
rect -6806 4837 -6803 4883
rect -6803 4837 -6757 4883
rect -6757 4837 -6754 4883
rect -6806 4834 -6754 4837
rect -6806 4763 -6754 4766
rect -6806 4717 -6803 4763
rect -6803 4717 -6757 4763
rect -6757 4717 -6754 4763
rect -6806 4714 -6754 4717
rect -7286 4283 -7234 4286
rect -7286 4237 -7283 4283
rect -7283 4237 -7237 4283
rect -7237 4237 -7234 4283
rect -7286 4234 -7234 4237
rect -6806 4043 -6754 4046
rect -6806 3997 -6803 4043
rect -6803 3997 -6757 4043
rect -6757 3997 -6754 4043
rect -6806 3994 -6754 3997
rect -6806 2843 -6754 2846
rect -6806 2797 -6803 2843
rect -6803 2797 -6757 2843
rect -6757 2797 -6754 2843
rect -6806 2794 -6754 2797
rect -6806 2363 -6754 2366
rect -6806 2317 -6803 2363
rect -6803 2317 -6757 2363
rect -6757 2317 -6754 2363
rect -6806 2314 -6754 2317
rect -6806 1883 -6754 1886
rect -6806 1837 -6803 1883
rect -6803 1837 -6757 1883
rect -6757 1837 -6754 1883
rect -6806 1834 -6754 1837
rect -6806 1403 -6754 1406
rect -6806 1357 -6803 1403
rect -6803 1357 -6757 1403
rect -6757 1357 -6754 1403
rect -6806 1354 -6754 1357
rect -6806 923 -6754 926
rect -6806 877 -6803 923
rect -6803 877 -6757 923
rect -6757 877 -6754 923
rect -6806 874 -6754 877
rect -6806 -277 -6754 -274
rect -6806 -323 -6803 -277
rect -6803 -323 -6757 -277
rect -6757 -323 -6754 -277
rect -6806 -326 -6754 -323
rect -6806 -757 -6754 -754
rect -6806 -803 -6803 -757
rect -6803 -803 -6757 -757
rect -6757 -803 -6754 -757
rect -6806 -806 -6754 -803
rect -6806 -877 -6754 -874
rect -6806 -923 -6803 -877
rect -6803 -923 -6757 -877
rect -6757 -923 -6754 -877
rect -6806 -926 -6754 -923
rect -6806 -997 -6754 -994
rect -6806 -1043 -6803 -997
rect -6803 -1043 -6757 -997
rect -6757 -1043 -6754 -997
rect -6806 -1046 -6754 -1043
rect -6806 -1237 -6754 -1234
rect -6806 -1283 -6803 -1237
rect -6803 -1283 -6757 -1237
rect -6757 -1283 -6754 -1237
rect -6806 -1286 -6754 -1283
<< metal2 >>
rect -6840 6808 -6720 6840
rect -6840 6752 -6808 6808
rect -6752 6752 -6720 6808
rect -6840 6568 -6720 6752
rect -6840 6512 -6808 6568
rect -6752 6512 -6720 6568
rect -6840 6448 -6720 6512
rect -6840 6392 -6808 6448
rect -6752 6392 -6720 6448
rect -6840 6328 -6720 6392
rect -6840 6272 -6808 6328
rect -6752 6272 -6720 6328
rect -6840 6240 -6720 6272
rect -7080 5848 -6960 5880
rect -7080 5792 -7048 5848
rect -6992 5792 -6960 5848
rect -7080 5368 -6960 5792
rect -7080 5312 -7048 5368
rect -6992 5312 -6960 5368
rect -7080 5280 -6960 5312
rect -6840 5368 -6720 5400
rect -6840 5312 -6808 5368
rect -6752 5312 -6720 5368
rect -6840 4886 -6720 5312
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4766 -6720 4834
rect -6840 4714 -6806 4766
rect -6754 4714 -6720 4766
rect -6840 4680 -6720 4714
rect -7320 4288 -7200 4320
rect -7320 4232 -7288 4288
rect -7232 4232 -7200 4288
rect -7320 4200 -7200 4232
rect -6840 4048 -6720 4080
rect -6840 3992 -6808 4048
rect -6752 3992 -6720 4048
rect -6840 2848 -6720 3992
rect -6840 2792 -6808 2848
rect -6752 2792 -6720 2848
rect -6840 2368 -6720 2792
rect -6840 2312 -6808 2368
rect -6752 2312 -6720 2368
rect -6840 1888 -6720 2312
rect -6840 1832 -6808 1888
rect -6752 1832 -6720 1888
rect -6840 1408 -6720 1832
rect -6840 1352 -6808 1408
rect -6752 1352 -6720 1408
rect -6840 928 -6720 1352
rect -6840 872 -6808 928
rect -6752 872 -6720 928
rect -6840 -272 -6720 872
rect -6840 -328 -6808 -272
rect -6752 -328 -6720 -272
rect -6840 -754 -6720 -328
rect -6840 -806 -6806 -754
rect -6754 -806 -6720 -754
rect -6840 -874 -6720 -806
rect -6840 -926 -6806 -874
rect -6754 -926 -6720 -874
rect -6840 -994 -6720 -926
rect -6840 -1046 -6806 -994
rect -6754 -1046 -6720 -994
rect -6840 -1232 -6720 -1046
rect -6840 -1288 -6808 -1232
rect -6752 -1288 -6720 -1232
rect -6840 -1320 -6720 -1288
<< via2 >>
rect -6808 6806 -6752 6808
rect -6808 6754 -6806 6806
rect -6806 6754 -6754 6806
rect -6754 6754 -6752 6806
rect -6808 6752 -6752 6754
rect -6808 6566 -6752 6568
rect -6808 6514 -6806 6566
rect -6806 6514 -6754 6566
rect -6754 6514 -6752 6566
rect -6808 6512 -6752 6514
rect -6808 6446 -6752 6448
rect -6808 6394 -6806 6446
rect -6806 6394 -6754 6446
rect -6754 6394 -6752 6446
rect -6808 6392 -6752 6394
rect -6808 6326 -6752 6328
rect -6808 6274 -6806 6326
rect -6806 6274 -6754 6326
rect -6754 6274 -6752 6326
rect -6808 6272 -6752 6274
rect -7048 5792 -6992 5848
rect -7048 5312 -6992 5368
rect -6808 5312 -6752 5368
rect -7288 4286 -7232 4288
rect -7288 4234 -7286 4286
rect -7286 4234 -7234 4286
rect -7234 4234 -7232 4286
rect -7288 4232 -7232 4234
rect -6808 4046 -6752 4048
rect -6808 3994 -6806 4046
rect -6806 3994 -6754 4046
rect -6754 3994 -6752 4046
rect -6808 3992 -6752 3994
rect -6808 2846 -6752 2848
rect -6808 2794 -6806 2846
rect -6806 2794 -6754 2846
rect -6754 2794 -6752 2846
rect -6808 2792 -6752 2794
rect -6808 2366 -6752 2368
rect -6808 2314 -6806 2366
rect -6806 2314 -6754 2366
rect -6754 2314 -6752 2366
rect -6808 2312 -6752 2314
rect -6808 1886 -6752 1888
rect -6808 1834 -6806 1886
rect -6806 1834 -6754 1886
rect -6754 1834 -6752 1886
rect -6808 1832 -6752 1834
rect -6808 1406 -6752 1408
rect -6808 1354 -6806 1406
rect -6806 1354 -6754 1406
rect -6754 1354 -6752 1406
rect -6808 1352 -6752 1354
rect -6808 926 -6752 928
rect -6808 874 -6806 926
rect -6806 874 -6754 926
rect -6754 874 -6752 926
rect -6808 872 -6752 874
rect -6808 -274 -6752 -272
rect -6808 -326 -6806 -274
rect -6806 -326 -6754 -274
rect -6754 -326 -6752 -274
rect -6808 -328 -6752 -326
rect -6808 -1234 -6752 -1232
rect -6808 -1286 -6806 -1234
rect -6806 -1286 -6754 -1234
rect -6754 -1286 -6752 -1234
rect -6808 -1288 -6752 -1286
<< metal3 >>
rect -7560 6808 -6600 6840
rect -7560 6752 -6808 6808
rect -6752 6752 -6600 6808
rect -7560 6568 -6600 6752
rect -7560 6512 -6808 6568
rect -6752 6512 -6600 6568
rect -7560 6448 -6600 6512
rect -7560 6392 -6808 6448
rect -6752 6392 -6600 6448
rect -7560 6328 -6600 6392
rect -7560 6272 -6808 6328
rect -6752 6272 -6600 6328
rect -7560 6240 -6600 6272
rect -7560 5848 -6600 5880
rect -7560 5792 -7048 5848
rect -6992 5792 -6600 5848
rect -7560 5700 -6600 5792
rect -7560 5520 -6600 5640
rect -7560 5368 -6600 5460
rect -7560 5312 -7048 5368
rect -6992 5312 -6808 5368
rect -6752 5312 -6600 5368
rect -7560 5280 -6600 5312
rect -7560 4288 -6600 4320
rect -7560 4232 -7288 4288
rect -7232 4232 -6600 4288
rect -7560 4200 -6600 4232
rect -7560 4048 -6600 4080
rect -7560 3992 -6808 4048
rect -6752 3992 -6600 4048
rect -7560 3960 -6600 3992
rect -7560 3540 -6600 3840
rect -7560 3360 -6600 3480
rect -7560 3000 -6600 3300
rect -7560 2848 -6600 2880
rect -7560 2792 -6808 2848
rect -6752 2792 -6600 2848
rect -7560 2760 -6600 2792
rect -7560 2520 -6600 2640
rect -7560 2368 -6600 2400
rect -7560 2312 -6808 2368
rect -6752 2312 -6600 2368
rect -7560 2280 -6600 2312
rect -7560 2040 -6600 2160
rect -7560 1888 -6600 1920
rect -7560 1832 -6808 1888
rect -6752 1832 -6600 1888
rect -7560 1800 -6600 1832
rect -7560 1560 -6600 1680
rect -7560 1408 -6600 1440
rect -7560 1352 -6808 1408
rect -6752 1352 -6600 1408
rect -7560 1320 -6600 1352
rect -7560 1080 -6600 1200
rect -7560 928 -6600 960
rect -7560 872 -6808 928
rect -6752 872 -6600 928
rect -7560 840 -6600 872
rect -7560 420 -6600 720
rect -7560 240 -6600 360
rect -7560 -120 -6600 180
rect -7560 -272 -6600 -240
rect -7560 -328 -6808 -272
rect -6752 -328 -6600 -272
rect -7560 -360 -6600 -328
rect -7560 -1232 -6600 -720
rect -7560 -1288 -6808 -1232
rect -6752 -1288 -6600 -1232
rect -7560 -1320 -6600 -1288
<< labels >>
rlabel metal1 s -7020 -540 -7020 -540 4 lo
rlabel metal1 s -7020 4500 -7020 4500 4 hi
rlabel metal1 s -7020 6060 -7020 6060 4 hih
rlabel metal3 s -7560 6240 -6600 6840 4 vdd
port 1 nsew
rlabel metal3 s -7560 5520 -6600 5640 4 gp
port 2 nsew
rlabel metal3 s -7560 4200 -6600 4320 4 bp
port 3 nsew
rlabel metal3 s -7560 5760 -6600 5880 4 vreg
port 4 nsew
rlabel metal3 s -7560 2520 -6600 2640 4 im
port 5 nsew
rlabel metal3 s -7560 1080 -6600 1200 4 ip
port 6 nsew
rlabel metal3 s -7560 -1320 -6600 -720 4 gnd
port 7 nsew
rlabel metal3 s -7560 3360 -6600 3480 4 xm
port 8 nsew
rlabel metal3 s -7560 3720 -6600 3840 4 op
port 9 nsew
rlabel metal3 s -7560 3000 -6600 3120 4 op
port 9 nsew
rlabel metal3 s -7560 240 -6600 360 4 xp
port 10 nsew
rlabel metal3 s -7560 -120 -6600 0 4 om
port 11 nsew
rlabel metal3 s -7560 600 -6600 720 4 om
port 11 nsew
rlabel metal3 s -7560 2040 -6600 2160 4 x
port 12 nsew
rlabel metal3 s -7560 1560 -6600 1680 4 y
port 13 nsew
<< end >>
