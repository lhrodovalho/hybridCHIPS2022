magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7380 5220 -6600 6420
rect -7380 3660 -6600 4980
<< nmos >>
rect -6960 -1080 -6840 -720
<< pmos >>
rect -6960 4200 -6840 4500
<< mvpmos >>
rect -6960 5760 -6840 6120
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
<< pdiff >>
rect -7080 4403 -6960 4500
rect -7080 4357 -7043 4403
rect -6997 4357 -6960 4403
rect -7080 4283 -6960 4357
rect -7080 4237 -7043 4283
rect -6997 4237 -6960 4283
rect -7080 4200 -6960 4237
rect -6840 4403 -6720 4500
rect -6840 4357 -6803 4403
rect -6757 4357 -6720 4403
rect -6840 4283 -6720 4357
rect -6840 4237 -6803 4283
rect -6757 4237 -6720 4283
rect -6840 4200 -6720 4237
<< mvpdiff >>
rect -7080 6083 -6960 6120
rect -7080 6037 -7043 6083
rect -6997 6037 -6960 6083
rect -7080 5963 -6960 6037
rect -7080 5917 -7043 5963
rect -6997 5917 -6960 5963
rect -7080 5843 -6960 5917
rect -7080 5797 -7043 5843
rect -6997 5797 -6960 5843
rect -7080 5760 -6960 5797
rect -6840 6083 -6720 6120
rect -6840 6037 -6803 6083
rect -6757 6037 -6720 6083
rect -6840 5963 -6720 6037
rect -6840 5917 -6803 5963
rect -6757 5917 -6720 5963
rect -6840 5843 -6720 5917
rect -6840 5797 -6803 5843
rect -6757 5797 -6720 5843
rect -6840 5760 -6720 5797
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
<< pdiffc >>
rect -7043 4357 -6997 4403
rect -7043 4237 -6997 4283
rect -6803 4357 -6757 4403
rect -6803 4237 -6757 4283
<< mvpdiffc >>
rect -7043 6037 -6997 6083
rect -7043 5917 -6997 5963
rect -7043 5797 -6997 5843
rect -6803 6037 -6757 6083
rect -6803 5917 -6757 5963
rect -6803 5797 -6757 5843
<< psubdiff >>
rect -7560 6563 -6600 6600
rect -7560 6517 -7523 6563
rect -7477 6517 -7403 6563
rect -7357 6517 -7283 6563
rect -7237 6517 -7163 6563
rect -7117 6517 -7043 6563
rect -6997 6517 -6923 6563
rect -6877 6517 -6803 6563
rect -6757 6517 -6683 6563
rect -6637 6517 -6600 6563
rect -7560 6480 -6600 6517
rect -7560 6443 -7440 6480
rect -7560 6397 -7523 6443
rect -7477 6397 -7440 6443
rect -7560 6323 -7440 6397
rect -7560 6277 -7523 6323
rect -7477 6277 -7440 6323
rect -7560 6203 -7440 6277
rect -7560 6157 -7523 6203
rect -7477 6157 -7440 6203
rect -7560 6083 -7440 6157
rect -7560 6037 -7523 6083
rect -7477 6037 -7440 6083
rect -7560 5963 -7440 6037
rect -7560 5917 -7523 5963
rect -7477 5917 -7440 5963
rect -7560 5843 -7440 5917
rect -7560 5797 -7523 5843
rect -7477 5797 -7440 5843
rect -7560 5723 -7440 5797
rect -7560 5677 -7523 5723
rect -7477 5677 -7440 5723
rect -7560 5603 -7440 5677
rect -7560 5557 -7523 5603
rect -7477 5557 -7440 5603
rect -7560 5483 -7440 5557
rect -7560 5437 -7523 5483
rect -7477 5437 -7440 5483
rect -7560 5363 -7440 5437
rect -7560 5317 -7523 5363
rect -7477 5317 -7440 5363
rect -7560 5243 -7440 5317
rect -7560 5197 -7523 5243
rect -7477 5197 -7440 5243
rect -7560 5160 -7440 5197
rect -7560 5123 -6600 5160
rect -7560 5077 -7523 5123
rect -7477 5077 -7403 5123
rect -7357 5077 -7283 5123
rect -7237 5077 -7163 5123
rect -7117 5077 -7043 5123
rect -6997 5077 -6923 5123
rect -6877 5077 -6803 5123
rect -6757 5077 -6683 5123
rect -6637 5077 -6600 5123
rect -7560 5040 -6600 5077
rect -7560 5003 -7440 5040
rect -7560 4957 -7523 5003
rect -7477 4957 -7440 5003
rect -7560 4883 -7440 4957
rect -7560 4837 -7523 4883
rect -7477 4837 -7440 4883
rect -7560 4763 -7440 4837
rect -7560 4717 -7523 4763
rect -7477 4717 -7440 4763
rect -7560 4643 -7440 4717
rect -7560 4597 -7523 4643
rect -7477 4597 -7440 4643
rect -7560 4523 -7440 4597
rect -7560 4477 -7523 4523
rect -7477 4477 -7440 4523
rect -7560 4403 -7440 4477
rect -7560 4357 -7523 4403
rect -7477 4357 -7440 4403
rect -7560 4283 -7440 4357
rect -7560 4237 -7523 4283
rect -7477 4237 -7440 4283
rect -7560 4163 -7440 4237
rect -7560 4117 -7523 4163
rect -7477 4117 -7440 4163
rect -7560 4043 -7440 4117
rect -7560 3997 -7523 4043
rect -7477 3997 -7440 4043
rect -7560 3923 -7440 3997
rect -7560 3877 -7523 3923
rect -7477 3877 -7440 3923
rect -7560 3803 -7440 3877
rect -7560 3757 -7523 3803
rect -7477 3757 -7440 3803
rect -7560 3683 -7440 3757
rect -7560 3637 -7523 3683
rect -7477 3637 -7440 3683
rect -7560 3600 -7440 3637
rect -7560 3563 -6600 3600
rect -7560 3517 -7523 3563
rect -7477 3517 -7403 3563
rect -7357 3517 -7283 3563
rect -7237 3517 -7163 3563
rect -7117 3517 -7043 3563
rect -6997 3517 -6923 3563
rect -6877 3517 -6803 3563
rect -6757 3517 -6683 3563
rect -6637 3517 -6600 3563
rect -7560 3480 -6600 3517
rect -7560 3443 -7440 3480
rect -7560 3397 -7523 3443
rect -7477 3397 -7440 3443
rect -7560 3323 -7440 3397
rect -7560 3277 -7523 3323
rect -7477 3277 -7440 3323
rect -7560 3203 -7440 3277
rect -7560 3157 -7523 3203
rect -7477 3157 -7440 3203
rect -7560 3083 -7440 3157
rect -7560 3037 -7523 3083
rect -7477 3037 -7440 3083
rect -7560 2963 -7440 3037
rect -7560 2917 -7523 2963
rect -7477 2917 -7440 2963
rect -7560 2843 -7440 2917
rect -7560 2797 -7523 2843
rect -7477 2797 -7440 2843
rect -7560 2723 -7440 2797
rect -7560 2677 -7523 2723
rect -7477 2677 -7440 2723
rect -7560 2640 -7440 2677
rect -7560 2603 -6600 2640
rect -7560 2557 -7523 2603
rect -7477 2557 -7403 2603
rect -7357 2557 -7283 2603
rect -7237 2557 -7163 2603
rect -7117 2557 -7043 2603
rect -6997 2557 -6923 2603
rect -6877 2557 -6803 2603
rect -6757 2557 -6683 2603
rect -6637 2557 -6600 2603
rect -7560 2520 -6600 2557
rect -7560 2483 -7440 2520
rect -7560 2437 -7523 2483
rect -7477 2437 -7440 2483
rect -7560 2363 -7440 2437
rect -7560 2317 -7523 2363
rect -7477 2317 -7440 2363
rect -7560 2243 -7440 2317
rect -7560 2197 -7523 2243
rect -7477 2197 -7440 2243
rect -7560 2160 -7440 2197
rect -7560 2123 -6600 2160
rect -7560 2077 -7523 2123
rect -7477 2077 -7403 2123
rect -7357 2077 -7283 2123
rect -7237 2077 -7163 2123
rect -7117 2077 -7043 2123
rect -6997 2077 -6923 2123
rect -6877 2077 -6803 2123
rect -6757 2077 -6683 2123
rect -6637 2077 -6600 2123
rect -7560 2040 -6600 2077
rect -7560 2003 -7440 2040
rect -7560 1957 -7523 2003
rect -7477 1957 -7440 2003
rect -7560 1883 -7440 1957
rect -7560 1837 -7523 1883
rect -7477 1837 -7440 1883
rect -7560 1763 -7440 1837
rect -7560 1717 -7523 1763
rect -7477 1717 -7440 1763
rect -7560 1680 -7440 1717
rect -7560 1643 -6600 1680
rect -7560 1597 -7523 1643
rect -7477 1597 -7403 1643
rect -7357 1597 -7283 1643
rect -7237 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6600 1643
rect -7560 1560 -6600 1597
rect -7560 1523 -7440 1560
rect -7560 1477 -7523 1523
rect -7477 1477 -7440 1523
rect -7560 1403 -7440 1477
rect -7560 1357 -7523 1403
rect -7477 1357 -7440 1403
rect -7560 1283 -7440 1357
rect -7560 1237 -7523 1283
rect -7477 1237 -7440 1283
rect -7560 1200 -7440 1237
rect -7560 1163 -6600 1200
rect -7560 1117 -7523 1163
rect -7477 1117 -7403 1163
rect -7357 1117 -7283 1163
rect -7237 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6600 1163
rect -7560 1080 -6600 1117
rect -7560 1043 -7440 1080
rect -7560 997 -7523 1043
rect -7477 997 -7440 1043
rect -7560 923 -7440 997
rect -7560 877 -7523 923
rect -7477 877 -7440 923
rect -7560 803 -7440 877
rect -7560 757 -7523 803
rect -7477 757 -7440 803
rect -7560 720 -7440 757
rect -7560 683 -6600 720
rect -7560 637 -7523 683
rect -7477 637 -7403 683
rect -7357 637 -7283 683
rect -7237 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6600 683
rect -7560 600 -6600 637
rect -7560 563 -7440 600
rect -7560 517 -7523 563
rect -7477 517 -7440 563
rect -7560 443 -7440 517
rect -7560 397 -7523 443
rect -7477 397 -7440 443
rect -7560 323 -7440 397
rect -7560 277 -7523 323
rect -7477 277 -7440 323
rect -7560 203 -7440 277
rect -7560 157 -7523 203
rect -7477 157 -7440 203
rect -7560 83 -7440 157
rect -7560 37 -7523 83
rect -7477 37 -7440 83
rect -7560 -37 -7440 37
rect -7560 -83 -7523 -37
rect -7477 -83 -7440 -37
rect -7560 -157 -7440 -83
rect -7560 -203 -7523 -157
rect -7477 -203 -7440 -157
rect -7560 -240 -7440 -203
rect -7560 -277 -6600 -240
rect -7560 -323 -7523 -277
rect -7477 -323 -7403 -277
rect -7357 -323 -7283 -277
rect -7237 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6600 -277
rect -7560 -360 -6600 -323
rect -7560 -397 -7440 -360
rect -7560 -443 -7523 -397
rect -7477 -443 -7440 -397
rect -7560 -517 -7440 -443
rect -7560 -563 -7523 -517
rect -7477 -563 -7440 -517
rect -7560 -637 -7440 -563
rect -7560 -683 -7523 -637
rect -7477 -683 -7440 -637
rect -7560 -757 -7440 -683
rect -7560 -803 -7523 -757
rect -7477 -803 -7440 -757
rect -7560 -877 -7440 -803
rect -7560 -923 -7523 -877
rect -7477 -923 -7440 -877
rect -7560 -997 -7440 -923
rect -7560 -1043 -7523 -997
rect -7477 -1043 -7440 -997
rect -7560 -1117 -7440 -1043
rect -7560 -1163 -7523 -1117
rect -7477 -1163 -7440 -1117
rect -7560 -1200 -7440 -1163
rect -7560 -1237 -6600 -1200
rect -7560 -1283 -7523 -1237
rect -7477 -1283 -7403 -1237
rect -7357 -1283 -7283 -1237
rect -7237 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6600 -1237
rect -7560 -1320 -6600 -1283
<< nsubdiff >>
rect -7320 4883 -6720 4920
rect -7320 4837 -7283 4883
rect -7237 4837 -7163 4883
rect -7117 4837 -7043 4883
rect -6997 4837 -6923 4883
rect -6877 4837 -6803 4883
rect -6757 4837 -6720 4883
rect -7320 4800 -6720 4837
rect -7320 4763 -7200 4800
rect -7320 4717 -7283 4763
rect -7237 4717 -7200 4763
rect -7320 4643 -7200 4717
rect -7320 4597 -7283 4643
rect -7237 4597 -7200 4643
rect -7320 4523 -7200 4597
rect -7320 4477 -7283 4523
rect -7237 4477 -7200 4523
rect -7320 4403 -7200 4477
rect -7320 4357 -7283 4403
rect -7237 4357 -7200 4403
rect -7320 4283 -7200 4357
rect -7320 4237 -7283 4283
rect -7237 4237 -7200 4283
rect -7320 4163 -7200 4237
rect -7320 4117 -7283 4163
rect -7237 4117 -7200 4163
rect -7320 4043 -7200 4117
rect -7320 3997 -7283 4043
rect -7237 3997 -7200 4043
rect -7320 3923 -7200 3997
rect -7320 3877 -7283 3923
rect -7237 3877 -7200 3923
rect -7320 3840 -7200 3877
rect -7320 3803 -6720 3840
rect -7320 3757 -7283 3803
rect -7237 3757 -7163 3803
rect -7117 3757 -7043 3803
rect -6997 3757 -6923 3803
rect -6877 3757 -6803 3803
rect -6757 3757 -6720 3803
rect -7320 3720 -6720 3757
<< mvnsubdiff >>
rect -7320 6323 -6720 6360
rect -7320 6277 -7283 6323
rect -7237 6277 -7163 6323
rect -7117 6277 -7043 6323
rect -6997 6277 -6923 6323
rect -6877 6277 -6803 6323
rect -6757 6277 -6720 6323
rect -7320 6240 -6720 6277
rect -7320 6203 -7200 6240
rect -7320 6157 -7283 6203
rect -7237 6157 -7200 6203
rect -7320 6083 -7200 6157
rect -7320 6037 -7283 6083
rect -7237 6037 -7200 6083
rect -7320 5963 -7200 6037
rect -7320 5917 -7283 5963
rect -7237 5917 -7200 5963
rect -7320 5843 -7200 5917
rect -7320 5797 -7283 5843
rect -7237 5797 -7200 5843
rect -7320 5723 -7200 5797
rect -7320 5677 -7283 5723
rect -7237 5677 -7200 5723
rect -7320 5603 -7200 5677
rect -7320 5557 -7283 5603
rect -7237 5557 -7200 5603
rect -7320 5483 -7200 5557
rect -7320 5437 -7283 5483
rect -7237 5437 -7200 5483
rect -7320 5400 -7200 5437
rect -7320 5363 -6720 5400
rect -7320 5317 -7283 5363
rect -7237 5317 -7163 5363
rect -7117 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6720 5363
rect -7320 5280 -6720 5317
<< psubdiffcont >>
rect -7523 6517 -7477 6563
rect -7403 6517 -7357 6563
rect -7283 6517 -7237 6563
rect -7163 6517 -7117 6563
rect -7043 6517 -6997 6563
rect -6923 6517 -6877 6563
rect -6803 6517 -6757 6563
rect -6683 6517 -6637 6563
rect -7523 6397 -7477 6443
rect -7523 6277 -7477 6323
rect -7523 6157 -7477 6203
rect -7523 6037 -7477 6083
rect -7523 5917 -7477 5963
rect -7523 5797 -7477 5843
rect -7523 5677 -7477 5723
rect -7523 5557 -7477 5603
rect -7523 5437 -7477 5483
rect -7523 5317 -7477 5363
rect -7523 5197 -7477 5243
rect -7523 5077 -7477 5123
rect -7403 5077 -7357 5123
rect -7283 5077 -7237 5123
rect -7163 5077 -7117 5123
rect -7043 5077 -6997 5123
rect -6923 5077 -6877 5123
rect -6803 5077 -6757 5123
rect -6683 5077 -6637 5123
rect -7523 4957 -7477 5003
rect -7523 4837 -7477 4883
rect -7523 4717 -7477 4763
rect -7523 4597 -7477 4643
rect -7523 4477 -7477 4523
rect -7523 4357 -7477 4403
rect -7523 4237 -7477 4283
rect -7523 4117 -7477 4163
rect -7523 3997 -7477 4043
rect -7523 3877 -7477 3923
rect -7523 3757 -7477 3803
rect -7523 3637 -7477 3683
rect -7523 3517 -7477 3563
rect -7403 3517 -7357 3563
rect -7283 3517 -7237 3563
rect -7163 3517 -7117 3563
rect -7043 3517 -6997 3563
rect -6923 3517 -6877 3563
rect -6803 3517 -6757 3563
rect -6683 3517 -6637 3563
rect -7523 3397 -7477 3443
rect -7523 3277 -7477 3323
rect -7523 3157 -7477 3203
rect -7523 3037 -7477 3083
rect -7523 2917 -7477 2963
rect -7523 2797 -7477 2843
rect -7523 2677 -7477 2723
rect -7523 2557 -7477 2603
rect -7403 2557 -7357 2603
rect -7283 2557 -7237 2603
rect -7163 2557 -7117 2603
rect -7043 2557 -6997 2603
rect -6923 2557 -6877 2603
rect -6803 2557 -6757 2603
rect -6683 2557 -6637 2603
rect -7523 2437 -7477 2483
rect -7523 2317 -7477 2363
rect -7523 2197 -7477 2243
rect -7523 2077 -7477 2123
rect -7403 2077 -7357 2123
rect -7283 2077 -7237 2123
rect -7163 2077 -7117 2123
rect -7043 2077 -6997 2123
rect -6923 2077 -6877 2123
rect -6803 2077 -6757 2123
rect -6683 2077 -6637 2123
rect -7523 1957 -7477 2003
rect -7523 1837 -7477 1883
rect -7523 1717 -7477 1763
rect -7523 1597 -7477 1643
rect -7403 1597 -7357 1643
rect -7283 1597 -7237 1643
rect -7163 1597 -7117 1643
rect -7043 1597 -6997 1643
rect -6923 1597 -6877 1643
rect -6803 1597 -6757 1643
rect -6683 1597 -6637 1643
rect -7523 1477 -7477 1523
rect -7523 1357 -7477 1403
rect -7523 1237 -7477 1283
rect -7523 1117 -7477 1163
rect -7403 1117 -7357 1163
rect -7283 1117 -7237 1163
rect -7163 1117 -7117 1163
rect -7043 1117 -6997 1163
rect -6923 1117 -6877 1163
rect -6803 1117 -6757 1163
rect -6683 1117 -6637 1163
rect -7523 997 -7477 1043
rect -7523 877 -7477 923
rect -7523 757 -7477 803
rect -7523 637 -7477 683
rect -7403 637 -7357 683
rect -7283 637 -7237 683
rect -7163 637 -7117 683
rect -7043 637 -6997 683
rect -6923 637 -6877 683
rect -6803 637 -6757 683
rect -6683 637 -6637 683
rect -7523 517 -7477 563
rect -7523 397 -7477 443
rect -7523 277 -7477 323
rect -7523 157 -7477 203
rect -7523 37 -7477 83
rect -7523 -83 -7477 -37
rect -7523 -203 -7477 -157
rect -7523 -323 -7477 -277
rect -7403 -323 -7357 -277
rect -7283 -323 -7237 -277
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -7523 -443 -7477 -397
rect -7523 -563 -7477 -517
rect -7523 -683 -7477 -637
rect -7523 -803 -7477 -757
rect -7523 -923 -7477 -877
rect -7523 -1043 -7477 -997
rect -7523 -1163 -7477 -1117
rect -7523 -1283 -7477 -1237
rect -7403 -1283 -7357 -1237
rect -7283 -1283 -7237 -1237
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
<< nsubdiffcont >>
rect -7283 4837 -7237 4883
rect -7163 4837 -7117 4883
rect -7043 4837 -6997 4883
rect -6923 4837 -6877 4883
rect -6803 4837 -6757 4883
rect -7283 4717 -7237 4763
rect -7283 4597 -7237 4643
rect -7283 4477 -7237 4523
rect -7283 4357 -7237 4403
rect -7283 4237 -7237 4283
rect -7283 4117 -7237 4163
rect -7283 3997 -7237 4043
rect -7283 3877 -7237 3923
rect -7283 3757 -7237 3803
rect -7163 3757 -7117 3803
rect -7043 3757 -6997 3803
rect -6923 3757 -6877 3803
rect -6803 3757 -6757 3803
<< mvnsubdiffcont >>
rect -7283 6277 -7237 6323
rect -7163 6277 -7117 6323
rect -7043 6277 -6997 6323
rect -6923 6277 -6877 6323
rect -6803 6277 -6757 6323
rect -7283 6157 -7237 6203
rect -7283 6037 -7237 6083
rect -7283 5917 -7237 5963
rect -7283 5797 -7237 5843
rect -7283 5677 -7237 5723
rect -7283 5557 -7237 5603
rect -7283 5437 -7237 5483
rect -7283 5317 -7237 5363
rect -7163 5317 -7117 5363
rect -7043 5317 -6997 5363
rect -6923 5317 -6877 5363
rect -6803 5317 -6757 5363
<< polysilicon >>
rect -6960 6120 -6840 6180
rect -6960 5603 -6840 5760
rect -6960 5557 -6923 5603
rect -6877 5557 -6840 5603
rect -6960 5520 -6840 5557
rect -6960 4500 -6840 4560
rect -6960 4043 -6840 4200
rect -6960 3997 -6923 4043
rect -6877 3997 -6840 4043
rect -6960 3960 -6840 3997
rect -6960 -517 -6840 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6840 -517
rect -6960 -720 -6840 -563
rect -6960 -1140 -6840 -1080
<< polycontact >>
rect -6923 5557 -6877 5603
rect -6923 3997 -6877 4043
rect -6923 -563 -6877 -517
<< metal1 >>
rect -7560 6563 -6600 6600
rect -7560 6517 -7523 6563
rect -7477 6517 -7403 6563
rect -7357 6517 -7283 6563
rect -7237 6517 -7163 6563
rect -7117 6517 -7043 6563
rect -6997 6517 -6923 6563
rect -6877 6517 -6803 6563
rect -6757 6517 -6683 6563
rect -6637 6517 -6600 6563
rect -7560 6480 -6600 6517
rect -7560 6443 -7440 6480
rect -7560 6397 -7523 6443
rect -7477 6397 -7440 6443
rect -7560 6323 -7440 6397
rect -7560 6277 -7523 6323
rect -7477 6277 -7440 6323
rect -7560 6203 -7440 6277
rect -7560 6157 -7523 6203
rect -7477 6157 -7440 6203
rect -7560 6083 -7440 6157
rect -7560 6037 -7523 6083
rect -7477 6037 -7440 6083
rect -7560 5963 -7440 6037
rect -7560 5917 -7523 5963
rect -7477 5917 -7440 5963
rect -7560 5843 -7440 5917
rect -7560 5797 -7523 5843
rect -7477 5797 -7440 5843
rect -7560 5723 -7440 5797
rect -7560 5677 -7523 5723
rect -7477 5677 -7440 5723
rect -7560 5603 -7440 5677
rect -7560 5557 -7523 5603
rect -7477 5557 -7440 5603
rect -7560 5483 -7440 5557
rect -7560 5437 -7523 5483
rect -7477 5437 -7440 5483
rect -7560 5363 -7440 5437
rect -7560 5317 -7523 5363
rect -7477 5317 -7440 5363
rect -7560 5243 -7440 5317
rect -7320 6326 -6600 6360
rect -7320 6323 -6806 6326
rect -7320 6277 -7283 6323
rect -7237 6277 -7163 6323
rect -7117 6277 -7043 6323
rect -6997 6277 -6923 6323
rect -6877 6277 -6806 6323
rect -7320 6274 -6806 6277
rect -6754 6274 -6600 6326
rect -7320 6240 -6600 6274
rect -7320 6203 -7200 6240
rect -7320 6157 -7283 6203
rect -7237 6157 -7200 6203
rect -7320 6083 -7200 6157
rect -7320 6037 -7283 6083
rect -7237 6037 -7200 6083
rect -7320 5963 -7200 6037
rect -7320 5917 -7283 5963
rect -7237 5917 -7200 5963
rect -7320 5843 -7200 5917
rect -7320 5797 -7283 5843
rect -7237 5797 -7200 5843
rect -7320 5723 -7200 5797
rect -7320 5677 -7283 5723
rect -7237 5677 -7200 5723
rect -7320 5603 -7200 5677
rect -7320 5557 -7283 5603
rect -7237 5557 -7200 5603
rect -7320 5483 -7200 5557
rect -7080 6083 -6960 6120
rect -7080 6037 -7043 6083
rect -6997 6037 -6960 6083
rect -7080 5963 -6960 6037
rect -7080 5917 -7043 5963
rect -6997 5917 -6960 5963
rect -7080 5843 -6960 5917
rect -7080 5797 -7043 5843
rect -6997 5797 -6960 5843
rect -7080 5640 -6960 5797
rect -6840 6086 -6720 6120
rect -6840 6034 -6806 6086
rect -6754 6034 -6720 6086
rect -6840 5966 -6720 6034
rect -6840 5914 -6806 5966
rect -6754 5914 -6720 5966
rect -6840 5846 -6720 5914
rect -6840 5794 -6806 5846
rect -6754 5794 -6720 5846
rect -6840 5760 -6720 5794
rect -7080 5603 -6840 5640
rect -7080 5557 -6923 5603
rect -6877 5557 -6840 5603
rect -7080 5520 -6840 5557
rect -7320 5437 -7283 5483
rect -7237 5437 -7200 5483
rect -7320 5400 -7200 5437
rect -7320 5363 -6600 5400
rect -7320 5317 -7283 5363
rect -7237 5317 -7163 5363
rect -7117 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6600 5363
rect -7320 5280 -6600 5317
rect -7560 5197 -7523 5243
rect -7477 5197 -7440 5243
rect -7560 5160 -7440 5197
rect -7560 5123 -6600 5160
rect -7560 5077 -7523 5123
rect -7477 5077 -7403 5123
rect -7357 5077 -7283 5123
rect -7237 5077 -7163 5123
rect -7117 5077 -7043 5123
rect -6997 5077 -6923 5123
rect -6877 5077 -6803 5123
rect -6757 5077 -6683 5123
rect -6637 5077 -6600 5123
rect -7560 5040 -6600 5077
rect -7560 5003 -7440 5040
rect -7560 4957 -7523 5003
rect -7477 4957 -7440 5003
rect -7560 4883 -7440 4957
rect -7560 4837 -7523 4883
rect -7477 4837 -7440 4883
rect -7560 4763 -7440 4837
rect -7560 4717 -7523 4763
rect -7477 4717 -7440 4763
rect -7560 4643 -7440 4717
rect -7560 4597 -7523 4643
rect -7477 4597 -7440 4643
rect -7560 4523 -7440 4597
rect -7560 4477 -7523 4523
rect -7477 4477 -7440 4523
rect -7560 4403 -7440 4477
rect -7560 4357 -7523 4403
rect -7477 4357 -7440 4403
rect -7560 4283 -7440 4357
rect -7560 4237 -7523 4283
rect -7477 4237 -7440 4283
rect -7560 4163 -7440 4237
rect -7560 4117 -7523 4163
rect -7477 4117 -7440 4163
rect -7560 4043 -7440 4117
rect -7560 3997 -7523 4043
rect -7477 3997 -7440 4043
rect -7560 3923 -7440 3997
rect -7560 3877 -7523 3923
rect -7477 3877 -7440 3923
rect -7560 3803 -7440 3877
rect -7560 3757 -7523 3803
rect -7477 3757 -7440 3803
rect -7560 3683 -7440 3757
rect -7320 4883 -6720 4920
rect -7320 4837 -7283 4883
rect -7237 4837 -7163 4883
rect -7117 4837 -7043 4883
rect -6997 4837 -6923 4883
rect -6877 4837 -6803 4883
rect -6757 4837 -6720 4883
rect -7320 4800 -6720 4837
rect -7320 4763 -7200 4800
rect -7320 4717 -7283 4763
rect -7237 4717 -7200 4763
rect -7320 4643 -7200 4717
rect -7320 4597 -7283 4643
rect -7237 4597 -7200 4643
rect -7320 4523 -7200 4597
rect -7320 4477 -7283 4523
rect -7237 4477 -7200 4523
rect -7320 4403 -7200 4477
rect -7320 4357 -7283 4403
rect -7237 4357 -7200 4403
rect -7320 4283 -7200 4357
rect -7320 4237 -7283 4283
rect -7237 4237 -7200 4283
rect -7320 4163 -7200 4237
rect -7320 4117 -7283 4163
rect -7237 4117 -7200 4163
rect -7320 4043 -7200 4117
rect -7320 3997 -7283 4043
rect -7237 3997 -7200 4043
rect -7320 3923 -7200 3997
rect -7080 4403 -6960 4500
rect -7080 4357 -7043 4403
rect -6997 4357 -6960 4403
rect -7080 4283 -6960 4357
rect -7080 4237 -7043 4283
rect -6997 4237 -6960 4283
rect -7080 4080 -6960 4237
rect -6840 4406 -6720 4500
rect -6840 4354 -6806 4406
rect -6754 4354 -6720 4406
rect -6840 4286 -6720 4354
rect -6840 4234 -6806 4286
rect -6754 4234 -6720 4286
rect -6840 4200 -6720 4234
rect -7080 4043 -6840 4080
rect -7080 3997 -6923 4043
rect -6877 3997 -6840 4043
rect -7080 3960 -6840 3997
rect -7320 3877 -7283 3923
rect -7237 3877 -7200 3923
rect -7320 3840 -7200 3877
rect -7320 3806 -6600 3840
rect -7320 3754 -7286 3806
rect -7234 3803 -6600 3806
rect -7234 3757 -7163 3803
rect -7117 3757 -7043 3803
rect -6997 3757 -6923 3803
rect -6877 3757 -6803 3803
rect -6757 3757 -6600 3803
rect -7234 3754 -6600 3757
rect -7320 3720 -6600 3754
rect -7560 3637 -7523 3683
rect -7477 3637 -7440 3683
rect -7560 3600 -7440 3637
rect -7560 3566 -6600 3600
rect -7560 3563 -6806 3566
rect -6754 3563 -6600 3566
rect -7560 3517 -7523 3563
rect -7477 3517 -7403 3563
rect -7357 3517 -7283 3563
rect -7237 3517 -7163 3563
rect -7117 3517 -7043 3563
rect -6997 3517 -6923 3563
rect -6877 3517 -6806 3563
rect -6754 3517 -6683 3563
rect -6637 3517 -6600 3563
rect -7560 3514 -6806 3517
rect -6754 3514 -6600 3517
rect -7560 3480 -6600 3514
rect -7560 3443 -7440 3480
rect -7560 3397 -7523 3443
rect -7477 3397 -7440 3443
rect -7560 3323 -7440 3397
rect -7560 3277 -7523 3323
rect -7477 3277 -7440 3323
rect -7560 3203 -7440 3277
rect -7560 3157 -7523 3203
rect -7477 3157 -7440 3203
rect -7560 3083 -7440 3157
rect -7560 3037 -7523 3083
rect -7477 3037 -7440 3083
rect -7560 2963 -7440 3037
rect -7560 2917 -7523 2963
rect -7477 2917 -7440 2963
rect -7560 2843 -7440 2917
rect -7560 2797 -7523 2843
rect -7477 2797 -7440 2843
rect -7560 2723 -7440 2797
rect -7560 2677 -7523 2723
rect -7477 2677 -7440 2723
rect -7560 2640 -7440 2677
rect -7560 2606 -6600 2640
rect -7560 2603 -6806 2606
rect -6754 2603 -6600 2606
rect -7560 2557 -7523 2603
rect -7477 2557 -7403 2603
rect -7357 2557 -7283 2603
rect -7237 2557 -7163 2603
rect -7117 2557 -7043 2603
rect -6997 2557 -6923 2603
rect -6877 2557 -6806 2603
rect -6754 2557 -6683 2603
rect -6637 2557 -6600 2603
rect -7560 2554 -6806 2557
rect -6754 2554 -6600 2557
rect -7560 2520 -6600 2554
rect -7560 2483 -7440 2520
rect -7560 2437 -7523 2483
rect -7477 2437 -7440 2483
rect -7560 2363 -7440 2437
rect -7560 2317 -7523 2363
rect -7477 2317 -7440 2363
rect -7560 2243 -7440 2317
rect -7560 2197 -7523 2243
rect -7477 2197 -7440 2243
rect -7560 2160 -7440 2197
rect -7560 2126 -6600 2160
rect -7560 2123 -6806 2126
rect -6754 2123 -6600 2126
rect -7560 2077 -7523 2123
rect -7477 2077 -7403 2123
rect -7357 2077 -7283 2123
rect -7237 2077 -7163 2123
rect -7117 2077 -7043 2123
rect -6997 2077 -6923 2123
rect -6877 2077 -6806 2123
rect -6754 2077 -6683 2123
rect -6637 2077 -6600 2123
rect -7560 2074 -6806 2077
rect -6754 2074 -6600 2077
rect -7560 2040 -6600 2074
rect -7560 2003 -7440 2040
rect -7560 1957 -7523 2003
rect -7477 1957 -7440 2003
rect -7560 1883 -7440 1957
rect -7560 1837 -7523 1883
rect -7477 1837 -7440 1883
rect -7560 1763 -7440 1837
rect -7560 1717 -7523 1763
rect -7477 1717 -7440 1763
rect -7560 1680 -7440 1717
rect -7560 1646 -6600 1680
rect -7560 1643 -6806 1646
rect -6754 1643 -6600 1646
rect -7560 1597 -7523 1643
rect -7477 1597 -7403 1643
rect -7357 1597 -7283 1643
rect -7237 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6806 1643
rect -6754 1597 -6683 1643
rect -6637 1597 -6600 1643
rect -7560 1594 -6806 1597
rect -6754 1594 -6600 1597
rect -7560 1560 -6600 1594
rect -7560 1523 -7440 1560
rect -7560 1477 -7523 1523
rect -7477 1477 -7440 1523
rect -7560 1403 -7440 1477
rect -7560 1357 -7523 1403
rect -7477 1357 -7440 1403
rect -7560 1283 -7440 1357
rect -7560 1237 -7523 1283
rect -7477 1237 -7440 1283
rect -7560 1200 -7440 1237
rect -7560 1166 -6600 1200
rect -7560 1163 -6806 1166
rect -6754 1163 -6600 1166
rect -7560 1117 -7523 1163
rect -7477 1117 -7403 1163
rect -7357 1117 -7283 1163
rect -7237 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6806 1163
rect -6754 1117 -6683 1163
rect -6637 1117 -6600 1163
rect -7560 1114 -6806 1117
rect -6754 1114 -6600 1117
rect -7560 1080 -6600 1114
rect -7560 1043 -7440 1080
rect -7560 997 -7523 1043
rect -7477 997 -7440 1043
rect -7560 923 -7440 997
rect -7560 877 -7523 923
rect -7477 877 -7440 923
rect -7560 803 -7440 877
rect -7560 757 -7523 803
rect -7477 757 -7440 803
rect -7560 720 -7440 757
rect -7560 686 -6600 720
rect -7560 683 -6806 686
rect -6754 683 -6600 686
rect -7560 637 -7523 683
rect -7477 637 -7403 683
rect -7357 637 -7283 683
rect -7237 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6806 683
rect -6754 637 -6683 683
rect -6637 637 -6600 683
rect -7560 634 -6806 637
rect -6754 634 -6600 637
rect -7560 600 -6600 634
rect -7560 563 -7440 600
rect -7560 517 -7523 563
rect -7477 517 -7440 563
rect -7560 443 -7440 517
rect -7560 397 -7523 443
rect -7477 397 -7440 443
rect -7560 323 -7440 397
rect -7560 277 -7523 323
rect -7477 277 -7440 323
rect -7560 203 -7440 277
rect -7560 157 -7523 203
rect -7477 157 -7440 203
rect -7560 83 -7440 157
rect -7560 37 -7523 83
rect -7477 37 -7440 83
rect -7560 -37 -7440 37
rect -7560 -83 -7523 -37
rect -7477 -83 -7440 -37
rect -7560 -157 -7440 -83
rect -7560 -203 -7523 -157
rect -7477 -203 -7440 -157
rect -7560 -240 -7440 -203
rect -7560 -274 -6600 -240
rect -7560 -277 -6806 -274
rect -6754 -277 -6600 -274
rect -7560 -323 -7523 -277
rect -7477 -323 -7403 -277
rect -7357 -323 -7283 -277
rect -7237 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6806 -277
rect -6754 -323 -6683 -277
rect -6637 -323 -6600 -277
rect -7560 -326 -6806 -323
rect -6754 -326 -6600 -323
rect -7560 -360 -6600 -326
rect -7560 -397 -7440 -360
rect -7560 -443 -7523 -397
rect -7477 -443 -7440 -397
rect -7560 -517 -7440 -443
rect -7560 -563 -7523 -517
rect -7477 -563 -7440 -517
rect -7560 -637 -7440 -563
rect -7560 -683 -7523 -637
rect -7477 -683 -7440 -637
rect -7560 -757 -7440 -683
rect -7560 -803 -7523 -757
rect -7477 -803 -7440 -757
rect -7560 -877 -7440 -803
rect -7560 -923 -7523 -877
rect -7477 -923 -7440 -877
rect -7560 -997 -7440 -923
rect -7560 -1043 -7523 -997
rect -7477 -1043 -7440 -997
rect -7560 -1117 -7440 -1043
rect -7080 -517 -6840 -480
rect -7080 -563 -6923 -517
rect -6877 -563 -6840 -517
rect -7080 -600 -6840 -563
rect -7080 -757 -6960 -600
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -754 -6720 -720
rect -6840 -806 -6806 -754
rect -6754 -806 -6720 -754
rect -6840 -874 -6720 -806
rect -6840 -926 -6806 -874
rect -6754 -926 -6720 -874
rect -6840 -994 -6720 -926
rect -6840 -1046 -6806 -994
rect -6754 -1046 -6720 -994
rect -6840 -1080 -6720 -1046
rect -7560 -1163 -7523 -1117
rect -7477 -1163 -7440 -1117
rect -7560 -1200 -7440 -1163
rect -7560 -1234 -6600 -1200
rect -7560 -1237 -6806 -1234
rect -6754 -1237 -6600 -1234
rect -7560 -1283 -7523 -1237
rect -7477 -1283 -7403 -1237
rect -7357 -1283 -7283 -1237
rect -7237 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6806 -1237
rect -6754 -1283 -6683 -1237
rect -6637 -1283 -6600 -1237
rect -7560 -1286 -6806 -1283
rect -6754 -1286 -6600 -1283
rect -7560 -1320 -6600 -1286
<< via1 >>
rect -6806 6323 -6754 6326
rect -6806 6277 -6803 6323
rect -6803 6277 -6757 6323
rect -6757 6277 -6754 6323
rect -6806 6274 -6754 6277
rect -6806 6083 -6754 6086
rect -6806 6037 -6803 6083
rect -6803 6037 -6757 6083
rect -6757 6037 -6754 6083
rect -6806 6034 -6754 6037
rect -6806 5963 -6754 5966
rect -6806 5917 -6803 5963
rect -6803 5917 -6757 5963
rect -6757 5917 -6754 5963
rect -6806 5914 -6754 5917
rect -6806 5843 -6754 5846
rect -6806 5797 -6803 5843
rect -6803 5797 -6757 5843
rect -6757 5797 -6754 5843
rect -6806 5794 -6754 5797
rect -6806 4403 -6754 4406
rect -6806 4357 -6803 4403
rect -6803 4357 -6757 4403
rect -6757 4357 -6754 4403
rect -6806 4354 -6754 4357
rect -6806 4283 -6754 4286
rect -6806 4237 -6803 4283
rect -6803 4237 -6757 4283
rect -6757 4237 -6754 4283
rect -6806 4234 -6754 4237
rect -7286 3803 -7234 3806
rect -7286 3757 -7283 3803
rect -7283 3757 -7237 3803
rect -7237 3757 -7234 3803
rect -7286 3754 -7234 3757
rect -6806 3563 -6754 3566
rect -6806 3517 -6803 3563
rect -6803 3517 -6757 3563
rect -6757 3517 -6754 3563
rect -6806 3514 -6754 3517
rect -6806 2603 -6754 2606
rect -6806 2557 -6803 2603
rect -6803 2557 -6757 2603
rect -6757 2557 -6754 2603
rect -6806 2554 -6754 2557
rect -6806 2123 -6754 2126
rect -6806 2077 -6803 2123
rect -6803 2077 -6757 2123
rect -6757 2077 -6754 2123
rect -6806 2074 -6754 2077
rect -6806 1643 -6754 1646
rect -6806 1597 -6803 1643
rect -6803 1597 -6757 1643
rect -6757 1597 -6754 1643
rect -6806 1594 -6754 1597
rect -6806 1163 -6754 1166
rect -6806 1117 -6803 1163
rect -6803 1117 -6757 1163
rect -6757 1117 -6754 1163
rect -6806 1114 -6754 1117
rect -6806 683 -6754 686
rect -6806 637 -6803 683
rect -6803 637 -6757 683
rect -6757 637 -6754 683
rect -6806 634 -6754 637
rect -6806 -277 -6754 -274
rect -6806 -323 -6803 -277
rect -6803 -323 -6757 -277
rect -6757 -323 -6754 -277
rect -6806 -326 -6754 -323
rect -6806 -757 -6754 -754
rect -6806 -803 -6803 -757
rect -6803 -803 -6757 -757
rect -6757 -803 -6754 -757
rect -6806 -806 -6754 -803
rect -6806 -877 -6754 -874
rect -6806 -923 -6803 -877
rect -6803 -923 -6757 -877
rect -6757 -923 -6754 -877
rect -6806 -926 -6754 -923
rect -6806 -997 -6754 -994
rect -6806 -1043 -6803 -997
rect -6803 -1043 -6757 -997
rect -6757 -1043 -6754 -997
rect -6806 -1046 -6754 -1043
rect -6806 -1237 -6754 -1234
rect -6806 -1283 -6803 -1237
rect -6803 -1283 -6757 -1237
rect -6757 -1283 -6754 -1237
rect -6806 -1286 -6754 -1283
<< metal2 >>
rect -6840 6328 -6720 6360
rect -6840 6272 -6808 6328
rect -6752 6272 -6720 6328
rect -6840 6088 -6720 6272
rect -6840 6032 -6808 6088
rect -6752 6032 -6720 6088
rect -6840 5968 -6720 6032
rect -6840 5912 -6808 5968
rect -6752 5912 -6720 5968
rect -6840 5848 -6720 5912
rect -6840 5792 -6808 5848
rect -6752 5792 -6720 5848
rect -6840 5760 -6720 5792
rect -7080 5368 -6960 5400
rect -7080 5312 -7048 5368
rect -6992 5312 -6960 5368
rect -7080 4888 -6960 5312
rect -7080 4832 -7048 4888
rect -6992 4832 -6960 4888
rect -7080 4800 -6960 4832
rect -6840 4888 -6720 4920
rect -6840 4832 -6808 4888
rect -6752 4832 -6720 4888
rect -6840 4406 -6720 4832
rect -6840 4354 -6806 4406
rect -6754 4354 -6720 4406
rect -6840 4286 -6720 4354
rect -6840 4234 -6806 4286
rect -6754 4234 -6720 4286
rect -6840 4200 -6720 4234
rect -7320 3808 -7200 3840
rect -7320 3752 -7288 3808
rect -7232 3752 -7200 3808
rect -7320 3720 -7200 3752
rect -6840 3568 -6720 3600
rect -6840 3512 -6808 3568
rect -6752 3512 -6720 3568
rect -6840 2608 -6720 3512
rect -6840 2552 -6808 2608
rect -6752 2552 -6720 2608
rect -6840 2128 -6720 2552
rect -6840 2072 -6808 2128
rect -6752 2072 -6720 2128
rect -6840 1648 -6720 2072
rect -6840 1592 -6808 1648
rect -6752 1592 -6720 1648
rect -6840 1168 -6720 1592
rect -6840 1112 -6808 1168
rect -6752 1112 -6720 1168
rect -6840 688 -6720 1112
rect -6840 632 -6808 688
rect -6752 632 -6720 688
rect -6840 -272 -6720 632
rect -6840 -328 -6808 -272
rect -6752 -328 -6720 -272
rect -6840 -754 -6720 -328
rect -6840 -806 -6806 -754
rect -6754 -806 -6720 -754
rect -6840 -874 -6720 -806
rect -6840 -926 -6806 -874
rect -6754 -926 -6720 -874
rect -6840 -994 -6720 -926
rect -6840 -1046 -6806 -994
rect -6754 -1046 -6720 -994
rect -6840 -1232 -6720 -1046
rect -6840 -1288 -6808 -1232
rect -6752 -1288 -6720 -1232
rect -6840 -1320 -6720 -1288
<< via2 >>
rect -6808 6326 -6752 6328
rect -6808 6274 -6806 6326
rect -6806 6274 -6754 6326
rect -6754 6274 -6752 6326
rect -6808 6272 -6752 6274
rect -6808 6086 -6752 6088
rect -6808 6034 -6806 6086
rect -6806 6034 -6754 6086
rect -6754 6034 -6752 6086
rect -6808 6032 -6752 6034
rect -6808 5966 -6752 5968
rect -6808 5914 -6806 5966
rect -6806 5914 -6754 5966
rect -6754 5914 -6752 5966
rect -6808 5912 -6752 5914
rect -6808 5846 -6752 5848
rect -6808 5794 -6806 5846
rect -6806 5794 -6754 5846
rect -6754 5794 -6752 5846
rect -6808 5792 -6752 5794
rect -7048 5312 -6992 5368
rect -7048 4832 -6992 4888
rect -6808 4832 -6752 4888
rect -7288 3806 -7232 3808
rect -7288 3754 -7286 3806
rect -7286 3754 -7234 3806
rect -7234 3754 -7232 3806
rect -7288 3752 -7232 3754
rect -6808 3566 -6752 3568
rect -6808 3514 -6806 3566
rect -6806 3514 -6754 3566
rect -6754 3514 -6752 3566
rect -6808 3512 -6752 3514
rect -6808 2606 -6752 2608
rect -6808 2554 -6806 2606
rect -6806 2554 -6754 2606
rect -6754 2554 -6752 2606
rect -6808 2552 -6752 2554
rect -6808 2126 -6752 2128
rect -6808 2074 -6806 2126
rect -6806 2074 -6754 2126
rect -6754 2074 -6752 2126
rect -6808 2072 -6752 2074
rect -6808 1646 -6752 1648
rect -6808 1594 -6806 1646
rect -6806 1594 -6754 1646
rect -6754 1594 -6752 1646
rect -6808 1592 -6752 1594
rect -6808 1166 -6752 1168
rect -6808 1114 -6806 1166
rect -6806 1114 -6754 1166
rect -6754 1114 -6752 1166
rect -6808 1112 -6752 1114
rect -6808 686 -6752 688
rect -6808 634 -6806 686
rect -6806 634 -6754 686
rect -6754 634 -6752 686
rect -6808 632 -6752 634
rect -6808 -274 -6752 -272
rect -6808 -326 -6806 -274
rect -6806 -326 -6754 -274
rect -6754 -326 -6752 -274
rect -6808 -328 -6752 -326
rect -6808 -1234 -6752 -1232
rect -6808 -1286 -6806 -1234
rect -6806 -1286 -6754 -1234
rect -6754 -1286 -6752 -1234
rect -6808 -1288 -6752 -1286
<< metal3 >>
rect -7560 6328 -6600 6360
rect -7560 6272 -6808 6328
rect -6752 6272 -6600 6328
rect -7560 6088 -6600 6272
rect -7560 6032 -6808 6088
rect -6752 6032 -6600 6088
rect -7560 5968 -6600 6032
rect -7560 5912 -6808 5968
rect -6752 5912 -6600 5968
rect -7560 5848 -6600 5912
rect -7560 5792 -6808 5848
rect -6752 5792 -6600 5848
rect -7560 5760 -6600 5792
rect -7560 5368 -6600 5400
rect -7560 5312 -7048 5368
rect -6992 5312 -6600 5368
rect -7560 5220 -6600 5312
rect -7560 5040 -6600 5160
rect -7560 4888 -6600 4980
rect -7560 4832 -7048 4888
rect -6992 4832 -6808 4888
rect -6752 4832 -6600 4888
rect -7560 4800 -6600 4832
rect -7560 3808 -6600 3840
rect -7560 3752 -7288 3808
rect -7232 3752 -6600 3808
rect -7560 3720 -6600 3752
rect -7560 3568 -6600 3600
rect -7560 3512 -6808 3568
rect -6752 3512 -6600 3568
rect -7560 3480 -6600 3512
rect -7560 2760 -6600 3360
rect -7560 2608 -6600 2640
rect -7560 2552 -6808 2608
rect -6752 2552 -6600 2608
rect -7560 2520 -6600 2552
rect -7560 2280 -6600 2400
rect -7560 2128 -6600 2160
rect -7560 2072 -6808 2128
rect -6752 2072 -6600 2128
rect -7560 2040 -6600 2072
rect -7560 1800 -6600 1920
rect -7560 1648 -6600 1680
rect -7560 1592 -6808 1648
rect -6752 1592 -6600 1648
rect -7560 1560 -6600 1592
rect -7560 1320 -6600 1440
rect -7560 1168 -6600 1200
rect -7560 1112 -6808 1168
rect -6752 1112 -6600 1168
rect -7560 1080 -6600 1112
rect -7560 840 -6600 960
rect -7560 688 -6600 720
rect -7560 632 -6808 688
rect -6752 632 -6600 688
rect -7560 600 -6600 632
rect -7560 -120 -6600 480
rect -7560 -272 -6600 -240
rect -7560 -328 -6808 -272
rect -6752 -328 -6600 -272
rect -7560 -360 -6600 -328
rect -7560 -1232 -6600 -720
rect -7560 -1288 -6808 -1232
rect -6752 -1288 -6600 -1232
rect -7560 -1320 -6600 -1288
<< labels >>
rlabel metal1 s -7020 5580 -7020 5580 4 hih
rlabel metal1 s -7020 4020 -7020 4020 4 hi
rlabel metal1 s -7020 -540 -7020 -540 4 lo
rlabel metal3 s -7560 5760 -6600 6360 4 vdd
port 1 nsew
rlabel metal3 s -7560 5280 -6600 5400 4 vreg
port 2 nsew
rlabel metal3 s -7560 5040 -6600 5160 4 gp
port 3 nsew
rlabel metal3 s -7560 3720 -6600 3840 4 bp
port 4 nsew
rlabel metal3 s -7560 2760 -6600 3360 4 op
port 5 nsew
rlabel metal3 s -7560 2280 -6600 2400 4 im
port 6 nsew
rlabel metal3 s -7560 1800 -6600 1920 4 x
port 7 nsew
rlabel metal3 s -7560 1320 -6600 1440 4 y
port 8 nsew
rlabel metal3 s -7560 840 -6600 960 4 ip
port 9 nsew
rlabel metal3 s -7560 -120 -6600 480 4 om
port 10 nsew
rlabel metal3 s -7560 -1320 -6600 -720 4 gnd
port 11 nsew
<< end >>
