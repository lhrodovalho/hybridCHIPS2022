* CMOS inverter-based single-ended amplifiers open-loop testbench

* Include GF180MCU device models
.include "../../../gf180mcuC/libs.tech/ngspice/design.ngspice"
.lib "../../../gf180mcuC/libs.tech/ngspice/sm141064.ngspice" statistical
.lib "../../../gf180mcuC/libs.tech/ngspice/sm141064.ngspice" mimcap_statistical
.temp 27

.param
+  sw_stat_global = 0
+  sw_stat_mismatch = 1

.include "../../inv/ngspice/inv.spice"
.include "../../nauta/magic/nauta.spice"
.include "../../barth/magic/barth.spice"
.include "../../manf/magic/manf.spice"
.include "../../barthmanf/magic/barthmanf.spice"
.include "../../barthnauta/magic/barthnauta.spice"
.include "../../nautanauta/magic/nautanauta.spice"
.include "../../nautavieru/magic/nautavieru.spice"
.include "../../manfvieru/magic/manfvieru.spice"

.param pVDD = 5.0
.param pC   = 10p
.param pIB  = 22u


VDD  vdd 0 dc {pVDD}
VSS  vss 0 0
ECM  cm vss vdd vss 0.5

vin in cm 0 ac 1
eip ip cm in cm -0.5
eim im cm in cm  0.5

vd0 vd0 vss dc {pVDD}
ib0 vdd ib0 {pIB}
xb0 ib0             vdd gp0 bp0 vreg0 vss inv_bias
x0  xp0 xm0 op0 om0 vd0 gp0 bp0 vreg0 vss nauta
cxp0 ip  xp0 1T
cxm0 im  xm0 1T
lop0 op0 xm0 1T
lom0 om0 xp0 1T
cop0 op0 cm  {pC}
com0 om0 cm  {pC}

vd1 vd1 vss dc {pVDD}
ib1 vdd ib1 {pIB}
xb1 ib1             vdd gp1 bp1 vreg1 vss inv_bias
x1  xp1 xm1 op1 om1 vd1 gp1 bp1 vreg1 vss barth
cxp1 ip  xp1 1T
cxm1 im  xm1 1T
lop1 op1 xm1 1T
lom1 om1 xp1 1T
cop1 op1 cm  {pC}
com1 om1 cm  {pC}

vd2 vd2 vss dc {pVDD}
ib2 vdd ib2 {pIB}
xb2 ib2             vdd gp2 bp2 vreg2 vss inv_bias
x2  xp2 xm2 op2 om2 vd2 gp2 bp2 vreg2 vss manf
cxp2 ip  xp2 1T
cxm2 im  xm2 1T
lop2 op2 xm2 1T
lom2 om2 xp2 1T
cop2 op2 cm  {pC}
com2 om2 cm  {pC}

vd3 vd3 vss dc {pVDD}
ib3 vdd ib3 {pIB}
xb3 ib3             vdd gp3 bp3 vreg3 vss inv_bias
x3  xp3 xm3 op3 om3 vd3 gp3 bp3 vreg3 vss barthnauta
cxp3 ip  xp3 1T
cxm3 im  xm3 1T
lop3 op3 xm3 1T
lom3 om3 xp3 1T
cop3 op3 cm  {pC}
com3 om3 cm  {pC}

vd4 vd4 vss dc {pVDD}
ib4 vdd ib4 {pIB}
xb4 ib4             vdd gp4 bp4 vreg4 vss inv_bias
x4  xp4 xm4 op4 om4 vd4 gp4 bp4 vreg4 vss barthmanf
cxp4 ip  xp4 1T
cxm4 im  xm4 1T
lop4 op4 xm4 1T
lom4 om4 xp4 1T
cop4 op4 cm  {pC}
com4 om4 cm  {pC}

vd5 vd5 vss dc {pVDD}
ib5 vdd ib5 {pIB}
xb5 ib5             vdd gp5 bp5 vreg5 vss inv_bias
x5  xp5 xm5 op5 om5 vd5 gp5 bp5 vreg5 vss nautanauta
cxp5 ip  xp5 1T
cxm5 im  xm5 1T
lop5 op5 xm5 1T
lom5 om5 xp5 1T
cop5 op5 cm  {pC}
com5 om5 cm  {pC}

vd6 vd6 vss dc {pVDD}
ib6 vdd ib6 {pIB}
xb6 ib6             vdd gp6 bp6 vreg6 vss inv_bias
x6  xp6 xm6 op6 om6 vd6 gp6 bp6 vreg6 vss nautavieru
cxp6 ip  xp6 1T
cxm6 im  xm6 1T
lop6 op6 xm6 1T
lom6 om6 xp6 1T
cop6 op6 cm  {pC}
com6 om6 cm  {pC}

vd7 vd7 vss dc {pVDD}
ib7 vdd ib7 {pIB}
xb7 ib7             vdd gp7 bp7 vreg7 vss inv_bias
x7  xp7 xm7 op7 om7 vd7 gp7 bp7 vreg7 vss manfvieru
cxp7 ip  xp7 1T
cxm7 im  xm7 1T
lop7 op7 xm7 1T
lom7 om7 xp7 1T
cop7 op7 cm  {pC}
com7 om7 cm  {pC}

.option gmin=1e-12

.control

	echo # Open-loop AC Monte Carlo simulation mismatch-only input voltage offset > ../data/ac_df_mc_mis_os.txt
	echo # N,B,M,BN,BM,NN,NV,MV >> ../data/ac_df_mc_mis_os.txt

	echo # Open-loop AC Monte Carlo simulation mismatch-only output common-voltage > ../data/ac_df_mc_mis_cm.txt
	echo # N,B,M,BN,BM,NN,NV,MV >> ../data/ac_df_mc_mis_cm.txt

	echo # Open-loop AC Monte Carlo simulation mismatch-only voltage gain > ../data/ac_df_mc_mis_av.txt
	echo # N,B,M,BN,BM,NN,NV,MV >> ../data/ac_df_mc_mis_av.txt

	echo # Open-loop AC Monte Carlo simulation mismatch-only GBW > ../data/ac_df_mc_mis_gbw.txt
	echo # N,B,M,BN,BM,NN,NV,MV >> ../data/ac_df_mc_mis_gbw.txt


	let run = 1
	dowhile run <= 100

	reset
	op

	let os0 = (op0-om0)
	let os1 = (op1-om1)
	let os2 = (op2-om2)
	let os3 = (op3-om3)
	let os4 = (op4-om4)
	let os5 = (op5-om5)
	let os6 = (op6-om6)
	let os7 = (op7-om7)

*	let cm0 = (op0+om7)/2
*	let cm1 = (op1+om7)/2
*	let cm2 = (op2+om7)/2
*	let cm3 = (op3+om7)/2
*	let cm4 = (op4+om7)/2
*	let cm5 = (op5+om7)/2
*	let cm6 = (op6+om7)/2
*	let cm7 = (op7+om7)/2

	let cm0 = (op0+om7-vreg0)/2
	let cm1 = (op1+om7-vreg1)/2
	let cm2 = (op2+om7-vreg2)/2
	let cm3 = (op3+om7-vreg3)/2
	let cm4 = (op4+om7-vreg4)/2
	let cm5 = (op5+om7-vreg5)/2
	let cm6 = (op6+om7-vreg6)/2
	let cm7 = (op7+om7-vreg7)/2

	let vreg0 = vreg0
	let vreg1 = vreg1
	let vreg2 = vreg2
	let vreg3 = vreg3
	let vreg4 = vreg4
	let vreg5 = vreg5
	let vreg6 = vreg6
	let vreg7 = vreg7

	echo $&os0,$&os1,$&os2,$&os3,$&os4,$&os5,$&os6,$&os7 >> ../data/ac_df_mc_mis_os.txt
	echo $&cm0,$&cm1,$&cm2,$&cm3,$&cm4,$&cm5,$&cm6,$&cm7 >> ../data/ac_df_mc_mis_cm.txt

	echo ">>> voltage offset"
	echo ">>> $&os0,$&os1,$&os2,$&os3,$&os4,$&os5,$&os6,$&os7"

	ac dec 100 1 1T

	let av0 = db(op0-om0)
	let av1 = db(op1-om1)
	let av2 = db(op2-om2)
	let av3 = db(op3-om3)
	let av4 = db(op4-om4)
	let av5 = db(op5-om5)
	let av6 = db(op6-om6)
	let av7 = db(op7-om7)
	
	let ph0 = cphase(op0-om0)*180/pi
	let ph1 = cphase(op1-om1)*180/pi
	let ph2 = cphase(op2-om2)*180/pi
	let ph3 = cphase(op3-om3)*180/pi
	let ph4 = cphase(op4-om4)*180/pi
	let ph5 = cphase(op5-om5)*180/pi
	let ph6 = cphase(op6-om6)*180/pi
	let ph7 = cphase(op7-om7)*180/pi

		
	meas ac gbw0 when av0=0
	meas ac gbw1 when av1=0
	meas ac gbw2 when av2=0
	meas ac gbw3 when av3=0
	meas ac gbw4 when av4=0
	meas ac gbw5 when av5=0
	meas ac gbw6 when av6=0
	meas ac gbw7 when av7=0
	
	meas ac pm0 find ph0 at=gbw0
	meas ac pm1 find ph1 at=gbw1
	meas ac pm2 find ph2 at=gbw2
	meas ac pm3 find ph3 at=gbw3
	meas ac pm4 find ph4 at=gbw4
	meas ac pm5 find ph5 at=gbw5
	meas ac pm6 find ph6 at=gbw6
	meas ac pm7 find ph7 at=gbw7
	
	meas ac av0_1khz find av0 at=1k
	meas ac av1_1khz find av1 at=1k
	meas ac av2_1khz find av2 at=1k
	meas ac av3_1khz find av3 at=1k
	meas ac av4_1khz find av4 at=1k
	meas ac av5_1khz find av5 at=1k
	meas ac av6_1khz find av6 at=1k
	meas ac av7_1khz find av7 at=1k
		
	echo $&av0_1khz,$&av1_1khz,$&av2_1khz,$&av3_1khz,$&av4_1khz,$&av5_1khz,$&av6_1khz,$&av7_1khz >> ../data/ac_df_mc_mis_av.txt
	echo $&gbw0,$&gbw1,$&gbw2,$&gbw3,$&gbw4,$&gbw5,$&gbw6,$&gbw7 >> ../data/ac_df_mc_mis_gbw.txt

	let run = run + 1
	end
		
.endc

.end
