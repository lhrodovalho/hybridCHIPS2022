magic
tech gf180mcuC
timestamp 1664012841
<< nwell >>
rect -720 522 -588 642
rect -720 366 -588 498
<< nmos >>
rect -696 -108 -684 -72
rect -672 -108 -660 -72
rect -648 -108 -636 -72
rect -624 -108 -612 -72
<< pmos >>
rect -696 420 -684 450
rect -672 420 -660 450
rect -648 420 -636 450
rect -624 420 -612 450
<< mvpmos >>
rect -696 576 -684 612
rect -672 576 -660 612
rect -648 576 -636 612
rect -624 576 -612 612
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
<< pdiff >>
rect -708 441 -696 450
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 429 -696 435
rect -708 423 -705 429
rect -699 423 -696 429
rect -708 420 -696 423
rect -684 441 -672 450
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 429 -672 435
rect -684 423 -681 429
rect -675 423 -672 429
rect -684 420 -672 423
rect -660 441 -648 450
rect -660 435 -657 441
rect -651 435 -648 441
rect -660 429 -648 435
rect -660 423 -657 429
rect -651 423 -648 429
rect -660 420 -648 423
rect -636 441 -624 450
rect -636 435 -633 441
rect -627 435 -624 441
rect -636 429 -624 435
rect -636 423 -633 429
rect -627 423 -624 429
rect -636 420 -624 423
rect -612 441 -600 450
rect -612 435 -609 441
rect -603 435 -600 441
rect -612 429 -600 435
rect -612 423 -609 429
rect -603 423 -600 429
rect -612 420 -600 423
<< mvpdiff >>
rect -708 609 -696 612
rect -708 603 -705 609
rect -699 603 -696 609
rect -708 597 -696 603
rect -708 591 -705 597
rect -699 591 -696 597
rect -708 585 -696 591
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 576 -696 579
rect -684 609 -672 612
rect -684 603 -681 609
rect -675 603 -672 609
rect -684 597 -672 603
rect -684 591 -681 597
rect -675 591 -672 597
rect -684 585 -672 591
rect -684 579 -681 585
rect -675 579 -672 585
rect -684 576 -672 579
rect -660 609 -648 612
rect -660 603 -657 609
rect -651 603 -648 609
rect -660 597 -648 603
rect -660 591 -657 597
rect -651 591 -648 597
rect -660 585 -648 591
rect -660 579 -657 585
rect -651 579 -648 585
rect -660 576 -648 579
rect -636 609 -624 612
rect -636 603 -633 609
rect -627 603 -624 609
rect -636 597 -624 603
rect -636 591 -633 597
rect -627 591 -624 597
rect -636 585 -624 591
rect -636 579 -633 585
rect -627 579 -624 585
rect -636 576 -624 579
rect -612 609 -600 612
rect -612 603 -609 609
rect -603 603 -600 609
rect -612 597 -600 603
rect -612 591 -609 597
rect -603 591 -600 597
rect -612 585 -600 591
rect -612 579 -609 585
rect -603 579 -600 585
rect -612 576 -600 579
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -633 -81 -627 -75
rect -633 -93 -627 -87
rect -633 -105 -627 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
<< pdiffc >>
rect -705 435 -699 441
rect -705 423 -699 429
rect -681 435 -675 441
rect -681 423 -675 429
rect -657 435 -651 441
rect -657 423 -651 429
rect -633 435 -627 441
rect -633 423 -627 429
rect -609 435 -603 441
rect -609 423 -603 429
<< mvpdiffc >>
rect -705 603 -699 609
rect -705 591 -699 597
rect -705 579 -699 585
rect -681 603 -675 609
rect -681 591 -675 597
rect -681 579 -675 585
rect -657 603 -651 609
rect -657 591 -651 597
rect -657 579 -651 585
rect -633 603 -627 609
rect -633 591 -627 597
rect -633 579 -627 585
rect -609 603 -603 609
rect -609 591 -603 597
rect -609 579 -603 585
<< psubdiff >>
rect -720 657 -588 660
rect -720 651 -717 657
rect -711 651 -705 657
rect -699 651 -693 657
rect -687 651 -681 657
rect -675 651 -669 657
rect -663 651 -657 657
rect -651 651 -645 657
rect -639 651 -633 657
rect -627 651 -621 657
rect -615 651 -609 657
rect -603 651 -597 657
rect -591 651 -588 657
rect -720 648 -588 651
rect -720 513 -588 516
rect -720 507 -717 513
rect -711 507 -705 513
rect -699 507 -693 513
rect -687 507 -681 513
rect -675 507 -669 513
rect -663 507 -657 513
rect -651 507 -645 513
rect -639 507 -633 513
rect -627 507 -621 513
rect -615 507 -609 513
rect -603 507 -597 513
rect -591 507 -588 513
rect -720 504 -588 507
rect -720 357 -588 360
rect -720 351 -717 357
rect -711 351 -705 357
rect -699 351 -693 357
rect -687 351 -681 357
rect -675 351 -669 357
rect -663 351 -657 357
rect -651 351 -645 357
rect -639 351 -633 357
rect -627 351 -621 357
rect -615 351 -609 357
rect -603 351 -597 357
rect -591 351 -588 357
rect -720 348 -588 351
rect -720 237 -588 240
rect -720 231 -717 237
rect -711 231 -705 237
rect -699 231 -693 237
rect -687 231 -681 237
rect -675 231 -669 237
rect -663 231 -657 237
rect -651 231 -645 237
rect -639 231 -633 237
rect -627 231 -621 237
rect -615 231 -609 237
rect -603 231 -597 237
rect -591 231 -588 237
rect -720 228 -588 231
rect -720 189 -588 192
rect -720 183 -717 189
rect -711 183 -705 189
rect -699 183 -693 189
rect -687 183 -681 189
rect -675 183 -669 189
rect -663 183 -657 189
rect -651 183 -645 189
rect -639 183 -633 189
rect -627 183 -621 189
rect -615 183 -609 189
rect -603 183 -597 189
rect -591 183 -588 189
rect -720 180 -588 183
rect -720 141 -588 144
rect -720 135 -717 141
rect -711 135 -705 141
rect -699 135 -693 141
rect -687 135 -681 141
rect -675 135 -669 141
rect -663 135 -657 141
rect -651 135 -645 141
rect -639 135 -633 141
rect -627 135 -621 141
rect -615 135 -609 141
rect -603 135 -597 141
rect -591 135 -588 141
rect -720 132 -588 135
rect -720 93 -588 96
rect -720 87 -717 93
rect -711 87 -705 93
rect -699 87 -693 93
rect -687 87 -681 93
rect -675 87 -669 93
rect -663 87 -657 93
rect -651 87 -645 93
rect -639 87 -633 93
rect -627 87 -621 93
rect -615 87 -609 93
rect -603 87 -597 93
rect -591 87 -588 93
rect -720 84 -588 87
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< nsubdiff >>
rect -708 489 -600 492
rect -708 483 -705 489
rect -699 483 -693 489
rect -687 483 -681 489
rect -675 483 -669 489
rect -663 483 -657 489
rect -651 483 -645 489
rect -639 483 -633 489
rect -627 483 -621 489
rect -615 483 -609 489
rect -603 483 -600 489
rect -708 480 -600 483
rect -708 381 -600 384
rect -708 375 -705 381
rect -699 375 -693 381
rect -687 375 -681 381
rect -675 375 -669 381
rect -663 375 -657 381
rect -651 375 -645 381
rect -639 375 -633 381
rect -627 375 -621 381
rect -615 375 -609 381
rect -603 375 -600 381
rect -708 372 -600 375
<< mvnsubdiff >>
rect -708 633 -600 636
rect -708 627 -705 633
rect -699 627 -693 633
rect -687 627 -681 633
rect -675 627 -669 633
rect -663 627 -657 633
rect -651 627 -645 633
rect -639 627 -633 633
rect -627 627 -621 633
rect -615 627 -609 633
rect -603 627 -600 633
rect -708 624 -600 627
rect -708 537 -600 540
rect -708 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -669 537
rect -663 531 -657 537
rect -651 531 -645 537
rect -639 531 -633 537
rect -627 531 -621 537
rect -615 531 -609 537
rect -603 531 -600 537
rect -708 528 -600 531
<< psubdiffcont >>
rect -717 651 -711 657
rect -705 651 -699 657
rect -693 651 -687 657
rect -681 651 -675 657
rect -669 651 -663 657
rect -657 651 -651 657
rect -645 651 -639 657
rect -633 651 -627 657
rect -621 651 -615 657
rect -609 651 -603 657
rect -597 651 -591 657
rect -717 507 -711 513
rect -705 507 -699 513
rect -693 507 -687 513
rect -681 507 -675 513
rect -669 507 -663 513
rect -657 507 -651 513
rect -645 507 -639 513
rect -633 507 -627 513
rect -621 507 -615 513
rect -609 507 -603 513
rect -597 507 -591 513
rect -717 351 -711 357
rect -705 351 -699 357
rect -693 351 -687 357
rect -681 351 -675 357
rect -669 351 -663 357
rect -657 351 -651 357
rect -645 351 -639 357
rect -633 351 -627 357
rect -621 351 -615 357
rect -609 351 -603 357
rect -597 351 -591 357
rect -717 231 -711 237
rect -705 231 -699 237
rect -693 231 -687 237
rect -681 231 -675 237
rect -669 231 -663 237
rect -657 231 -651 237
rect -645 231 -639 237
rect -633 231 -627 237
rect -621 231 -615 237
rect -609 231 -603 237
rect -597 231 -591 237
rect -717 183 -711 189
rect -705 183 -699 189
rect -693 183 -687 189
rect -681 183 -675 189
rect -669 183 -663 189
rect -657 183 -651 189
rect -645 183 -639 189
rect -633 183 -627 189
rect -621 183 -615 189
rect -609 183 -603 189
rect -597 183 -591 189
rect -717 135 -711 141
rect -705 135 -699 141
rect -693 135 -687 141
rect -681 135 -675 141
rect -669 135 -663 141
rect -657 135 -651 141
rect -645 135 -639 141
rect -633 135 -627 141
rect -621 135 -615 141
rect -609 135 -603 141
rect -597 135 -591 141
rect -717 87 -711 93
rect -705 87 -699 93
rect -693 87 -687 93
rect -681 87 -675 93
rect -669 87 -663 93
rect -657 87 -651 93
rect -645 87 -639 93
rect -633 87 -627 93
rect -621 87 -615 93
rect -609 87 -603 93
rect -597 87 -591 93
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -657 -33 -651 -27
rect -645 -33 -639 -27
rect -633 -33 -627 -27
rect -621 -33 -615 -27
rect -609 -33 -603 -27
rect -597 -33 -591 -27
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
rect -657 -129 -651 -123
rect -645 -129 -639 -123
rect -633 -129 -627 -123
rect -621 -129 -615 -123
rect -609 -129 -603 -123
rect -597 -129 -591 -123
<< nsubdiffcont >>
rect -705 483 -699 489
rect -693 483 -687 489
rect -681 483 -675 489
rect -669 483 -663 489
rect -657 483 -651 489
rect -645 483 -639 489
rect -633 483 -627 489
rect -621 483 -615 489
rect -609 483 -603 489
rect -705 375 -699 381
rect -693 375 -687 381
rect -681 375 -675 381
rect -669 375 -663 381
rect -657 375 -651 381
rect -645 375 -639 381
rect -633 375 -627 381
rect -621 375 -615 381
rect -609 375 -603 381
<< mvnsubdiffcont >>
rect -705 627 -699 633
rect -693 627 -687 633
rect -681 627 -675 633
rect -669 627 -663 633
rect -657 627 -651 633
rect -645 627 -639 633
rect -633 627 -627 633
rect -621 627 -615 633
rect -609 627 -603 633
rect -705 531 -699 537
rect -693 531 -687 537
rect -681 531 -675 537
rect -669 531 -663 537
rect -657 531 -651 537
rect -645 531 -639 537
rect -633 531 -627 537
rect -621 531 -615 537
rect -609 531 -603 537
<< polysilicon >>
rect -696 612 -684 618
rect -672 612 -660 618
rect -648 612 -636 618
rect -624 612 -612 618
rect -696 564 -684 576
rect -672 564 -660 576
rect -648 564 -636 576
rect -624 564 -612 576
rect -696 561 -612 564
rect -696 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -657 561
rect -651 555 -645 561
rect -639 555 -633 561
rect -627 555 -621 561
rect -615 555 -612 561
rect -696 552 -612 555
rect -696 450 -684 456
rect -672 450 -660 456
rect -648 450 -636 456
rect -624 450 -612 456
rect -696 408 -684 420
rect -672 408 -660 420
rect -696 405 -660 408
rect -696 399 -693 405
rect -687 399 -681 405
rect -675 399 -669 405
rect -663 399 -660 405
rect -696 396 -660 399
rect -648 408 -636 420
rect -624 408 -612 420
rect -648 405 -612 408
rect -648 399 -645 405
rect -639 399 -633 405
rect -627 399 -621 405
rect -615 399 -612 405
rect -648 396 -612 399
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -696 -72 -684 -60
rect -672 -72 -660 -60
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -648 -72 -636 -60
rect -624 -72 -612 -60
rect -696 -114 -684 -108
rect -672 -114 -660 -108
rect -648 -114 -636 -108
rect -624 -114 -612 -108
<< polycontact >>
rect -693 555 -687 561
rect -681 555 -675 561
rect -669 555 -663 561
rect -657 555 -651 561
rect -645 555 -639 561
rect -633 555 -627 561
rect -621 555 -615 561
rect -693 399 -687 405
rect -681 399 -675 405
rect -669 399 -663 405
rect -645 399 -639 405
rect -633 399 -627 405
rect -621 399 -615 405
rect -693 -57 -687 -51
rect -681 -57 -675 -51
rect -669 -57 -663 -51
rect -645 -57 -639 -51
rect -633 -57 -627 -51
rect -621 -57 -615 -51
<< metal1 >>
rect -720 657 -588 660
rect -720 651 -717 657
rect -711 651 -705 657
rect -699 651 -693 657
rect -687 651 -681 657
rect -675 651 -669 657
rect -663 651 -657 657
rect -651 651 -645 657
rect -639 651 -633 657
rect -627 651 -621 657
rect -615 651 -609 657
rect -603 651 -597 657
rect -591 651 -588 657
rect -720 648 -588 651
rect -720 633 -588 636
rect -720 627 -705 633
rect -699 627 -693 633
rect -687 627 -681 633
rect -675 627 -669 633
rect -663 627 -657 633
rect -651 627 -645 633
rect -639 627 -633 633
rect -627 627 -621 633
rect -615 627 -609 633
rect -603 627 -588 633
rect -720 624 -588 627
rect -708 609 -696 612
rect -708 603 -705 609
rect -699 603 -696 609
rect -708 597 -696 603
rect -708 591 -705 597
rect -699 591 -696 597
rect -708 585 -696 591
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 576 -696 579
rect -684 609 -672 612
rect -684 603 -681 609
rect -675 603 -672 609
rect -684 597 -672 603
rect -684 591 -681 597
rect -675 591 -672 597
rect -684 585 -672 591
rect -684 579 -681 585
rect -675 579 -672 585
rect -684 576 -672 579
rect -660 609 -648 612
rect -660 603 -657 609
rect -651 603 -648 609
rect -660 597 -648 603
rect -660 591 -657 597
rect -651 591 -648 597
rect -660 585 -648 591
rect -660 579 -657 585
rect -651 579 -648 585
rect -660 576 -648 579
rect -636 609 -624 612
rect -636 603 -633 609
rect -627 603 -624 609
rect -636 597 -624 603
rect -636 591 -633 597
rect -627 591 -624 597
rect -636 585 -624 591
rect -636 579 -633 585
rect -627 579 -624 585
rect -636 576 -624 579
rect -612 609 -600 612
rect -612 603 -609 609
rect -603 603 -600 609
rect -612 597 -600 603
rect -612 591 -609 597
rect -603 591 -600 597
rect -612 585 -600 591
rect -612 579 -609 585
rect -603 579 -600 585
rect -612 576 -600 579
rect -696 561 -612 564
rect -696 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -657 561
rect -651 555 -645 561
rect -639 555 -633 561
rect -627 555 -621 561
rect -615 555 -612 561
rect -696 552 -612 555
rect -720 537 -588 540
rect -720 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -669 537
rect -663 531 -657 537
rect -651 531 -645 537
rect -639 531 -633 537
rect -627 531 -621 537
rect -615 531 -609 537
rect -603 531 -588 537
rect -720 528 -588 531
rect -720 513 -588 516
rect -720 507 -717 513
rect -711 507 -705 513
rect -699 507 -693 513
rect -687 507 -681 513
rect -675 507 -669 513
rect -663 507 -657 513
rect -651 507 -645 513
rect -639 507 -633 513
rect -627 507 -621 513
rect -615 507 -609 513
rect -603 507 -597 513
rect -591 507 -588 513
rect -720 504 -588 507
rect -720 489 -588 492
rect -720 483 -705 489
rect -699 483 -693 489
rect -687 483 -681 489
rect -675 483 -669 489
rect -663 483 -657 489
rect -651 483 -645 489
rect -639 483 -633 489
rect -627 483 -621 489
rect -615 483 -609 489
rect -603 483 -588 489
rect -720 480 -588 483
rect -708 465 -600 468
rect -708 459 -705 465
rect -699 459 -657 465
rect -651 459 -609 465
rect -603 459 -600 465
rect -708 456 -600 459
rect -708 453 -696 456
rect -708 447 -705 453
rect -699 447 -696 453
rect -660 453 -648 456
rect -708 441 -696 447
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 429 -696 435
rect -708 423 -705 429
rect -699 423 -696 429
rect -708 420 -696 423
rect -684 441 -672 450
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 429 -672 435
rect -684 423 -681 429
rect -675 423 -672 429
rect -684 420 -672 423
rect -660 447 -657 453
rect -651 447 -648 453
rect -612 453 -600 456
rect -660 441 -648 447
rect -660 435 -657 441
rect -651 435 -648 441
rect -660 429 -648 435
rect -660 423 -657 429
rect -651 423 -648 429
rect -660 420 -648 423
rect -636 441 -624 450
rect -636 435 -633 441
rect -627 435 -624 441
rect -636 429 -624 435
rect -636 423 -633 429
rect -627 423 -624 429
rect -636 420 -624 423
rect -612 447 -609 453
rect -603 447 -600 453
rect -612 441 -600 447
rect -612 435 -609 441
rect -603 435 -600 441
rect -612 429 -600 435
rect -612 423 -609 429
rect -603 423 -600 429
rect -612 420 -600 423
rect -696 405 -660 408
rect -696 399 -693 405
rect -687 399 -681 405
rect -675 399 -669 405
rect -663 399 -660 405
rect -696 396 -660 399
rect -648 405 -612 408
rect -648 399 -645 405
rect -639 399 -633 405
rect -627 399 -621 405
rect -615 399 -612 405
rect -648 396 -612 399
rect -720 381 -588 384
rect -720 375 -705 381
rect -699 375 -693 381
rect -687 375 -681 381
rect -675 375 -669 381
rect -663 375 -657 381
rect -651 375 -645 381
rect -639 375 -633 381
rect -627 375 -621 381
rect -615 375 -609 381
rect -603 375 -588 381
rect -720 372 -588 375
rect -720 357 -588 360
rect -720 351 -717 357
rect -711 351 -705 357
rect -699 351 -693 357
rect -687 351 -681 357
rect -675 351 -669 357
rect -663 351 -657 357
rect -651 351 -645 357
rect -639 351 -633 357
rect -627 351 -621 357
rect -615 351 -609 357
rect -603 351 -597 357
rect -591 351 -588 357
rect -720 348 -588 351
rect -720 237 -588 240
rect -720 231 -717 237
rect -711 231 -705 237
rect -699 231 -693 237
rect -687 231 -681 237
rect -675 231 -669 237
rect -663 231 -657 237
rect -651 231 -645 237
rect -639 231 -633 237
rect -627 231 -621 237
rect -615 231 -609 237
rect -603 231 -597 237
rect -591 231 -588 237
rect -720 228 -588 231
rect -720 189 -588 192
rect -720 183 -717 189
rect -711 183 -705 189
rect -699 183 -693 189
rect -687 183 -681 189
rect -675 183 -669 189
rect -663 183 -657 189
rect -651 183 -645 189
rect -639 183 -633 189
rect -627 183 -621 189
rect -615 183 -609 189
rect -603 183 -597 189
rect -591 183 -588 189
rect -720 180 -588 183
rect -720 141 -588 144
rect -720 135 -717 141
rect -711 135 -705 141
rect -699 135 -693 141
rect -687 135 -681 141
rect -675 135 -669 141
rect -663 135 -657 141
rect -651 135 -645 141
rect -639 135 -633 141
rect -627 135 -621 141
rect -615 135 -609 141
rect -603 135 -597 141
rect -591 135 -588 141
rect -720 132 -588 135
rect -720 93 -588 96
rect -720 87 -717 93
rect -711 87 -705 93
rect -699 87 -693 93
rect -687 87 -681 93
rect -675 87 -669 93
rect -663 87 -657 93
rect -651 87 -645 93
rect -639 87 -633 93
rect -627 87 -621 93
rect -615 87 -609 93
rect -603 87 -597 93
rect -591 87 -588 93
rect -720 84 -588 87
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< via1 >>
rect -705 627 -699 633
rect -657 627 -651 633
rect -609 627 -603 633
rect -705 603 -699 609
rect -705 591 -699 597
rect -705 579 -699 585
rect -681 603 -675 609
rect -681 591 -675 597
rect -681 579 -675 585
rect -657 603 -651 609
rect -657 591 -651 597
rect -657 579 -651 585
rect -633 603 -627 609
rect -633 591 -627 597
rect -633 579 -627 585
rect -609 603 -603 609
rect -609 591 -603 597
rect -609 579 -603 585
rect -657 555 -651 561
rect -705 459 -699 465
rect -657 459 -651 465
rect -609 459 -603 465
rect -705 447 -699 453
rect -705 435 -699 441
rect -705 423 -699 429
rect -681 435 -675 441
rect -681 423 -675 429
rect -657 447 -651 453
rect -633 435 -627 441
rect -633 423 -627 429
rect -609 447 -603 453
rect -609 435 -603 441
rect -609 423 -603 429
rect -681 399 -675 405
rect -633 399 -627 405
rect -705 375 -699 381
rect -609 375 -603 381
rect -705 351 -699 357
rect -609 351 -603 357
rect -705 231 -699 237
rect -609 231 -603 237
rect -705 183 -699 189
rect -609 183 -603 189
rect -705 135 -699 141
rect -609 135 -603 141
rect -705 87 -699 93
rect -609 87 -603 93
rect -705 -33 -699 -27
rect -609 -33 -603 -27
rect -681 -57 -675 -51
rect -633 -57 -627 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal2 >>
rect -708 633 -696 636
rect -708 627 -705 633
rect -699 627 -696 633
rect -708 609 -696 627
rect -660 633 -648 636
rect -660 627 -657 633
rect -651 627 -648 633
rect -708 603 -705 609
rect -699 603 -696 609
rect -708 597 -696 603
rect -708 591 -705 597
rect -699 591 -696 597
rect -708 585 -696 591
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 576 -696 579
rect -684 609 -672 612
rect -684 603 -681 609
rect -675 603 -672 609
rect -684 597 -672 603
rect -684 591 -681 597
rect -675 591 -672 597
rect -684 585 -672 591
rect -684 579 -681 585
rect -675 579 -672 585
rect -684 537 -672 579
rect -660 609 -648 627
rect -612 633 -600 636
rect -612 627 -609 633
rect -603 627 -600 633
rect -660 603 -657 609
rect -651 603 -648 609
rect -660 597 -648 603
rect -660 591 -657 597
rect -651 591 -648 597
rect -660 585 -648 591
rect -660 579 -657 585
rect -651 579 -648 585
rect -660 576 -648 579
rect -636 609 -624 612
rect -636 603 -633 609
rect -627 603 -624 609
rect -636 597 -624 603
rect -636 591 -633 597
rect -627 591 -624 597
rect -636 585 -624 591
rect -636 579 -633 585
rect -627 579 -624 585
rect -660 561 -648 564
rect -660 555 -657 561
rect -651 555 -648 561
rect -660 552 -648 555
rect -684 531 -681 537
rect -675 531 -672 537
rect -708 489 -696 492
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 465 -696 483
rect -684 489 -672 531
rect -636 537 -624 579
rect -612 609 -600 627
rect -612 603 -609 609
rect -603 603 -600 609
rect -612 597 -600 603
rect -612 591 -609 597
rect -603 591 -600 597
rect -612 585 -600 591
rect -612 579 -609 585
rect -603 579 -600 585
rect -612 576 -600 579
rect -636 531 -633 537
rect -627 531 -624 537
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -660 489 -648 492
rect -660 483 -657 489
rect -651 483 -648 489
rect -708 459 -705 465
rect -699 459 -696 465
rect -708 453 -696 459
rect -708 447 -705 453
rect -699 447 -696 453
rect -660 465 -648 483
rect -636 489 -624 531
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 480 -624 483
rect -612 489 -600 492
rect -612 483 -609 489
rect -603 483 -600 489
rect -660 459 -657 465
rect -651 459 -648 465
rect -660 453 -648 459
rect -708 441 -696 447
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 429 -696 435
rect -708 423 -705 429
rect -699 423 -696 429
rect -708 420 -696 423
rect -684 441 -672 450
rect -660 447 -657 453
rect -651 447 -648 453
rect -612 465 -600 483
rect -612 459 -609 465
rect -603 459 -600 465
rect -612 453 -600 459
rect -660 444 -648 447
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 432 -672 435
rect -636 441 -624 450
rect -636 435 -633 441
rect -627 435 -624 441
rect -636 432 -624 435
rect -684 429 -624 432
rect -684 423 -681 429
rect -675 423 -633 429
rect -627 423 -624 429
rect -684 420 -624 423
rect -612 447 -609 453
rect -603 447 -600 453
rect -612 441 -600 447
rect -612 435 -609 441
rect -603 435 -600 441
rect -612 429 -600 435
rect -612 423 -609 429
rect -603 423 -600 429
rect -612 420 -600 423
rect -684 405 -672 408
rect -684 399 -681 405
rect -675 399 -672 405
rect -684 396 -672 399
rect -708 381 -696 384
rect -708 375 -705 381
rect -699 375 -696 381
rect -708 372 -696 375
rect -708 357 -696 360
rect -708 351 -705 357
rect -699 351 -696 357
rect -708 237 -696 351
rect -708 231 -705 237
rect -699 231 -696 237
rect -708 189 -696 231
rect -708 183 -705 189
rect -699 183 -696 189
rect -708 141 -696 183
rect -708 135 -705 141
rect -699 135 -696 141
rect -708 93 -696 135
rect -708 87 -705 93
rect -699 87 -696 93
rect -708 -27 -696 87
rect -708 -33 -705 -27
rect -699 -33 -696 -27
rect -708 -75 -696 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -123 -696 -105
rect -660 -75 -648 420
rect -636 405 -624 408
rect -636 399 -633 405
rect -627 399 -624 405
rect -636 396 -624 399
rect -612 381 -600 384
rect -612 375 -609 381
rect -603 375 -600 381
rect -612 372 -600 375
rect -612 357 -600 360
rect -612 351 -609 357
rect -603 351 -600 357
rect -612 237 -600 351
rect -612 231 -609 237
rect -603 231 -600 237
rect -612 189 -600 231
rect -612 183 -609 189
rect -603 183 -600 189
rect -612 141 -600 183
rect -612 135 -609 141
rect -603 135 -600 141
rect -612 93 -600 135
rect -612 87 -609 93
rect -603 87 -600 93
rect -612 -27 -600 87
rect -612 -33 -609 -27
rect -603 -33 -600 -27
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -612 -75 -600 -33
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -708 -129 -705 -123
rect -699 -129 -696 -123
rect -708 -132 -696 -129
rect -612 -123 -600 -105
rect -612 -129 -609 -123
rect -603 -129 -600 -123
rect -612 -132 -600 -129
<< via2 >>
rect -705 627 -699 633
rect -657 627 -651 633
rect -705 603 -699 609
rect -705 591 -699 597
rect -705 579 -699 585
rect -609 627 -603 633
rect -657 603 -651 609
rect -657 591 -651 597
rect -657 579 -651 585
rect -657 555 -651 561
rect -681 531 -675 537
rect -705 483 -699 489
rect -609 603 -603 609
rect -609 591 -603 597
rect -609 579 -603 585
rect -633 531 -627 537
rect -681 483 -675 489
rect -657 483 -651 489
rect -633 483 -627 489
rect -609 483 -603 489
rect -681 399 -675 405
rect -705 375 -699 381
rect -705 351 -699 357
rect -705 231 -699 237
rect -705 183 -699 189
rect -705 135 -699 141
rect -705 87 -699 93
rect -705 -33 -699 -27
rect -681 -57 -675 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -633 399 -627 405
rect -609 375 -603 381
rect -609 351 -603 357
rect -609 231 -603 237
rect -609 183 -603 189
rect -609 135 -603 141
rect -609 87 -603 93
rect -609 -33 -603 -27
rect -633 -57 -627 -51
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal3 >>
rect -720 633 -588 636
rect -720 627 -705 633
rect -699 627 -657 633
rect -651 627 -609 633
rect -603 627 -588 633
rect -720 609 -588 627
rect -720 603 -705 609
rect -699 603 -657 609
rect -651 603 -609 609
rect -603 603 -588 609
rect -720 597 -588 603
rect -720 591 -705 597
rect -699 591 -657 597
rect -651 591 -609 597
rect -603 591 -588 597
rect -720 585 -588 591
rect -720 579 -705 585
rect -699 579 -657 585
rect -651 579 -609 585
rect -603 579 -588 585
rect -720 576 -588 579
rect -660 561 -648 564
rect -660 555 -657 561
rect -651 555 -648 561
rect -660 552 -648 555
rect -720 537 -588 540
rect -720 531 -681 537
rect -675 531 -633 537
rect -627 531 -588 537
rect -720 522 -588 531
rect -720 513 -588 516
rect -720 507 -657 513
rect -651 507 -588 513
rect -720 504 -588 507
rect -720 489 -588 498
rect -720 483 -705 489
rect -699 483 -681 489
rect -675 483 -657 489
rect -651 483 -633 489
rect -627 483 -609 489
rect -603 483 -588 489
rect -720 480 -588 483
rect -684 405 -672 408
rect -684 399 -681 405
rect -675 399 -672 405
rect -684 396 -672 399
rect -636 405 -624 408
rect -636 399 -633 405
rect -627 399 -624 405
rect -636 396 -624 399
rect -720 381 -588 384
rect -720 375 -705 381
rect -699 375 -609 381
rect -603 375 -588 381
rect -720 372 -588 375
rect -720 357 -588 360
rect -720 351 -705 357
rect -699 351 -609 357
rect -603 351 -588 357
rect -720 348 -588 351
rect -720 306 -588 336
rect -720 288 -588 300
rect -720 252 -588 282
rect -720 237 -588 240
rect -720 231 -705 237
rect -699 231 -609 237
rect -603 231 -588 237
rect -720 228 -588 231
rect -720 204 -588 216
rect -720 189 -588 192
rect -720 183 -705 189
rect -699 183 -609 189
rect -603 183 -588 189
rect -720 180 -588 183
rect -720 156 -588 168
rect -720 141 -588 144
rect -720 135 -705 141
rect -699 135 -609 141
rect -603 135 -588 141
rect -720 132 -588 135
rect -720 108 -588 120
rect -720 93 -588 96
rect -720 87 -705 93
rect -699 87 -609 93
rect -603 87 -588 93
rect -720 84 -588 87
rect -720 42 -588 72
rect -720 24 -588 36
rect -720 -12 -588 18
rect -720 -27 -588 -24
rect -720 -33 -705 -27
rect -699 -33 -609 -27
rect -603 -33 -588 -27
rect -720 -36 -588 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -720 -75 -588 -72
rect -720 -81 -705 -75
rect -699 -81 -609 -75
rect -603 -81 -588 -75
rect -720 -87 -588 -81
rect -720 -93 -705 -87
rect -699 -93 -609 -87
rect -603 -93 -588 -87
rect -720 -99 -588 -93
rect -720 -105 -705 -99
rect -699 -105 -609 -99
rect -603 -105 -588 -99
rect -720 -123 -588 -105
rect -720 -129 -705 -123
rect -699 -129 -609 -123
rect -603 -129 -588 -123
rect -720 -132 -588 -129
<< via3 >>
rect -657 555 -651 561
rect -681 531 -675 537
rect -633 531 -627 537
rect -657 507 -651 513
rect -705 483 -699 489
rect -681 483 -675 489
rect -633 483 -627 489
rect -609 483 -603 489
rect -681 399 -675 405
rect -633 399 -627 405
rect -681 -57 -675 -51
rect -633 -57 -627 -51
<< metal4 >>
rect -660 561 -648 564
rect -660 555 -657 561
rect -651 555 -648 561
rect -684 537 -672 540
rect -684 531 -681 537
rect -675 531 -672 537
rect -708 489 -696 492
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 480 -696 483
rect -684 489 -672 531
rect -660 513 -648 555
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 504 -648 507
rect -636 537 -624 540
rect -636 531 -633 537
rect -627 531 -624 537
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -636 489 -624 531
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 480 -624 483
rect -612 489 -600 492
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 480 -600 483
rect -684 405 -672 408
rect -684 399 -681 405
rect -675 399 -672 405
rect -684 384 -672 399
rect -708 372 -672 384
rect -684 -51 -672 372
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 405 -624 408
rect -636 399 -633 405
rect -627 399 -624 405
rect -636 384 -624 399
rect -636 372 -600 384
rect -636 -51 -624 372
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
<< labels >>
rlabel metal4 -684 -12 -672 240 0 inl
port 1 nsew
rlabel metal4 -636 -12 -624 240 0 inr
port 2 nsew
rlabel metal2 -660 -12 -648 240 0 out
port 3 nsew
rlabel metal3 -720 -132 -588 -72 0 gnd
port 14 nsew
rlabel metal1 -684 -108 -672 -72 0 dl
rlabel metal1 -636 -108 -624 -72 0 dr
rlabel metal3 -720 -12 -588 0 0 om
port 15 nsew
rlabel metal3 -720 24 -588 36 0 xp
port 13 nsew
rlabel metal3 -720 108 -588 120 0 ip
port 11 nsew
rlabel metal3 -720 60 -588 72 0 om
port 15 nsew
rlabel metal3 -720 204 -588 216 0 im
port 10 nsew
rlabel metal3 -720 288 -588 300 0 xm
port 9 nsew
rlabel metal3 -720 576 -588 636 0 vdd
port 4 nsew
rlabel metal3 -720 504 -708 516 0 gp
port 5 nsew
rlabel metal3 -720 372 -708 384 0 bp
port 6 nsew
rlabel metal3 -720 528 -708 540 0 vreg
port 7 nsew
rlabel metal3 -720 324 -588 336 0 op
port 8 nsew
rlabel metal1 -708 504 -696 516 0 gnd
rlabel metal1 -708 648 -696 660 0 gnd
rlabel metal3 -720 252 -588 264 0 op
port 8 nsew
rlabel metal3 -720 156 -588 168 0 x
port 16 nsew
<< end >>
