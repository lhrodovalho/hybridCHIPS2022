magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7200 4260 -5880 5460
rect -7200 2700 -5880 4020
<< nmos >>
rect -6960 -1080 -6840 -720
rect -6720 -1080 -6600 -720
rect -6480 -1080 -6360 -720
rect -6240 -1080 -6120 -720
<< pmos >>
rect -6960 3240 -6840 3540
rect -6720 3240 -6600 3540
rect -6480 3240 -6360 3540
rect -6240 3240 -6120 3540
<< mvpmos >>
rect -6960 4800 -6840 5160
rect -6720 4800 -6600 5160
rect -6480 4800 -6360 5160
rect -6240 4800 -6120 5160
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -757 -6480 -720
rect -6600 -803 -6563 -757
rect -6517 -803 -6480 -757
rect -6600 -877 -6480 -803
rect -6600 -923 -6563 -877
rect -6517 -923 -6480 -877
rect -6600 -997 -6480 -923
rect -6600 -1043 -6563 -997
rect -6517 -1043 -6480 -997
rect -6600 -1080 -6480 -1043
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -757 -6000 -720
rect -6120 -803 -6083 -757
rect -6037 -803 -6000 -757
rect -6120 -877 -6000 -803
rect -6120 -923 -6083 -877
rect -6037 -923 -6000 -877
rect -6120 -997 -6000 -923
rect -6120 -1043 -6083 -997
rect -6037 -1043 -6000 -997
rect -6120 -1080 -6000 -1043
<< pdiff >>
rect -7080 3443 -6960 3540
rect -7080 3397 -7043 3443
rect -6997 3397 -6960 3443
rect -7080 3323 -6960 3397
rect -7080 3277 -7043 3323
rect -6997 3277 -6960 3323
rect -7080 3240 -6960 3277
rect -6840 3443 -6720 3540
rect -6840 3397 -6803 3443
rect -6757 3397 -6720 3443
rect -6840 3323 -6720 3397
rect -6840 3277 -6803 3323
rect -6757 3277 -6720 3323
rect -6840 3240 -6720 3277
rect -6600 3443 -6480 3540
rect -6600 3397 -6563 3443
rect -6517 3397 -6480 3443
rect -6600 3323 -6480 3397
rect -6600 3277 -6563 3323
rect -6517 3277 -6480 3323
rect -6600 3240 -6480 3277
rect -6360 3443 -6240 3540
rect -6360 3397 -6323 3443
rect -6277 3397 -6240 3443
rect -6360 3323 -6240 3397
rect -6360 3277 -6323 3323
rect -6277 3277 -6240 3323
rect -6360 3240 -6240 3277
rect -6120 3443 -6000 3540
rect -6120 3397 -6083 3443
rect -6037 3397 -6000 3443
rect -6120 3323 -6000 3397
rect -6120 3277 -6083 3323
rect -6037 3277 -6000 3323
rect -6120 3240 -6000 3277
<< mvpdiff >>
rect -7080 5123 -6960 5160
rect -7080 5077 -7043 5123
rect -6997 5077 -6960 5123
rect -7080 5003 -6960 5077
rect -7080 4957 -7043 5003
rect -6997 4957 -6960 5003
rect -7080 4883 -6960 4957
rect -7080 4837 -7043 4883
rect -6997 4837 -6960 4883
rect -7080 4800 -6960 4837
rect -6840 5123 -6720 5160
rect -6840 5077 -6803 5123
rect -6757 5077 -6720 5123
rect -6840 5003 -6720 5077
rect -6840 4957 -6803 5003
rect -6757 4957 -6720 5003
rect -6840 4883 -6720 4957
rect -6840 4837 -6803 4883
rect -6757 4837 -6720 4883
rect -6840 4800 -6720 4837
rect -6600 5123 -6480 5160
rect -6600 5077 -6563 5123
rect -6517 5077 -6480 5123
rect -6600 5003 -6480 5077
rect -6600 4957 -6563 5003
rect -6517 4957 -6480 5003
rect -6600 4883 -6480 4957
rect -6600 4837 -6563 4883
rect -6517 4837 -6480 4883
rect -6600 4800 -6480 4837
rect -6360 5123 -6240 5160
rect -6360 5077 -6323 5123
rect -6277 5077 -6240 5123
rect -6360 5003 -6240 5077
rect -6360 4957 -6323 5003
rect -6277 4957 -6240 5003
rect -6360 4883 -6240 4957
rect -6360 4837 -6323 4883
rect -6277 4837 -6240 4883
rect -6360 4800 -6240 4837
rect -6120 5123 -6000 5160
rect -6120 5077 -6083 5123
rect -6037 5077 -6000 5123
rect -6120 5003 -6000 5077
rect -6120 4957 -6083 5003
rect -6037 4957 -6000 5003
rect -6120 4883 -6000 4957
rect -6120 4837 -6083 4883
rect -6037 4837 -6000 4883
rect -6120 4800 -6000 4837
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
rect -6563 -803 -6517 -757
rect -6563 -923 -6517 -877
rect -6563 -1043 -6517 -997
rect -6323 -803 -6277 -757
rect -6323 -923 -6277 -877
rect -6323 -1043 -6277 -997
rect -6083 -803 -6037 -757
rect -6083 -923 -6037 -877
rect -6083 -1043 -6037 -997
<< pdiffc >>
rect -7043 3397 -6997 3443
rect -7043 3277 -6997 3323
rect -6803 3397 -6757 3443
rect -6803 3277 -6757 3323
rect -6563 3397 -6517 3443
rect -6563 3277 -6517 3323
rect -6323 3397 -6277 3443
rect -6323 3277 -6277 3323
rect -6083 3397 -6037 3443
rect -6083 3277 -6037 3323
<< mvpdiffc >>
rect -7043 5077 -6997 5123
rect -7043 4957 -6997 5003
rect -7043 4837 -6997 4883
rect -6803 5077 -6757 5123
rect -6803 4957 -6757 5003
rect -6803 4837 -6757 4883
rect -6563 5077 -6517 5123
rect -6563 4957 -6517 5003
rect -6563 4837 -6517 4883
rect -6323 5077 -6277 5123
rect -6323 4957 -6277 5003
rect -6323 4837 -6277 4883
rect -6083 5077 -6037 5123
rect -6083 4957 -6037 5003
rect -6083 4837 -6037 4883
<< psubdiff >>
rect -7200 5603 -5880 5640
rect -7200 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6563 5603
rect -6517 5557 -6443 5603
rect -6397 5557 -6323 5603
rect -6277 5557 -6203 5603
rect -6157 5557 -6083 5603
rect -6037 5557 -5963 5603
rect -5917 5557 -5880 5603
rect -7200 5520 -5880 5557
rect -7200 4163 -5880 4200
rect -7200 4117 -7163 4163
rect -7117 4117 -7043 4163
rect -6997 4117 -6923 4163
rect -6877 4117 -6803 4163
rect -6757 4117 -6683 4163
rect -6637 4117 -6563 4163
rect -6517 4117 -6443 4163
rect -6397 4117 -6323 4163
rect -6277 4117 -6203 4163
rect -6157 4117 -6083 4163
rect -6037 4117 -5963 4163
rect -5917 4117 -5880 4163
rect -7200 4080 -5880 4117
rect -7200 2603 -5880 2640
rect -7200 2557 -7163 2603
rect -7117 2557 -7043 2603
rect -6997 2557 -6923 2603
rect -6877 2557 -6803 2603
rect -6757 2557 -6683 2603
rect -6637 2557 -6563 2603
rect -6517 2557 -6443 2603
rect -6397 2557 -6323 2603
rect -6277 2557 -6203 2603
rect -6157 2557 -6083 2603
rect -6037 2557 -5963 2603
rect -5917 2557 -5880 2603
rect -7200 2520 -5880 2557
rect -7200 1643 -5880 1680
rect -7200 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6563 1643
rect -6517 1597 -6443 1643
rect -6397 1597 -6323 1643
rect -6277 1597 -6203 1643
rect -6157 1597 -6083 1643
rect -6037 1597 -5963 1643
rect -5917 1597 -5880 1643
rect -7200 1560 -5880 1597
rect -7200 1163 -5880 1200
rect -7200 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6563 1163
rect -6517 1117 -6443 1163
rect -6397 1117 -6323 1163
rect -6277 1117 -6203 1163
rect -6157 1117 -6083 1163
rect -6037 1117 -5963 1163
rect -5917 1117 -5880 1163
rect -7200 1080 -5880 1117
rect -7200 683 -5880 720
rect -7200 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6563 683
rect -6517 637 -6443 683
rect -6397 637 -6323 683
rect -6277 637 -6203 683
rect -6157 637 -6083 683
rect -6037 637 -5963 683
rect -5917 637 -5880 683
rect -7200 600 -5880 637
rect -7200 -277 -5880 -240
rect -7200 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6083 -277
rect -6037 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -360 -5880 -323
rect -7200 -1237 -5880 -1200
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6083 -1237
rect -6037 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1320 -5880 -1283
<< nsubdiff >>
rect -7080 3923 -6000 3960
rect -7080 3877 -7043 3923
rect -6997 3877 -6923 3923
rect -6877 3877 -6803 3923
rect -6757 3877 -6683 3923
rect -6637 3877 -6563 3923
rect -6517 3877 -6443 3923
rect -6397 3877 -6323 3923
rect -6277 3877 -6203 3923
rect -6157 3877 -6083 3923
rect -6037 3877 -6000 3923
rect -7080 3840 -6000 3877
rect -7080 2843 -6000 2880
rect -7080 2797 -7043 2843
rect -6997 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6683 2843
rect -6637 2797 -6563 2843
rect -6517 2797 -6443 2843
rect -6397 2797 -6323 2843
rect -6277 2797 -6203 2843
rect -6157 2797 -6083 2843
rect -6037 2797 -6000 2843
rect -7080 2760 -6000 2797
<< mvnsubdiff >>
rect -7080 5363 -6000 5400
rect -7080 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6683 5363
rect -6637 5317 -6563 5363
rect -6517 5317 -6443 5363
rect -6397 5317 -6323 5363
rect -6277 5317 -6203 5363
rect -6157 5317 -6083 5363
rect -6037 5317 -6000 5363
rect -7080 5280 -6000 5317
rect -7080 4403 -6000 4440
rect -7080 4357 -7043 4403
rect -6997 4357 -6923 4403
rect -6877 4357 -6803 4403
rect -6757 4357 -6683 4403
rect -6637 4357 -6563 4403
rect -6517 4357 -6443 4403
rect -6397 4357 -6323 4403
rect -6277 4357 -6203 4403
rect -6157 4357 -6083 4403
rect -6037 4357 -6000 4403
rect -7080 4320 -6000 4357
<< psubdiffcont >>
rect -7163 5557 -7117 5603
rect -7043 5557 -6997 5603
rect -6923 5557 -6877 5603
rect -6803 5557 -6757 5603
rect -6683 5557 -6637 5603
rect -6563 5557 -6517 5603
rect -6443 5557 -6397 5603
rect -6323 5557 -6277 5603
rect -6203 5557 -6157 5603
rect -6083 5557 -6037 5603
rect -5963 5557 -5917 5603
rect -7163 4117 -7117 4163
rect -7043 4117 -6997 4163
rect -6923 4117 -6877 4163
rect -6803 4117 -6757 4163
rect -6683 4117 -6637 4163
rect -6563 4117 -6517 4163
rect -6443 4117 -6397 4163
rect -6323 4117 -6277 4163
rect -6203 4117 -6157 4163
rect -6083 4117 -6037 4163
rect -5963 4117 -5917 4163
rect -7163 2557 -7117 2603
rect -7043 2557 -6997 2603
rect -6923 2557 -6877 2603
rect -6803 2557 -6757 2603
rect -6683 2557 -6637 2603
rect -6563 2557 -6517 2603
rect -6443 2557 -6397 2603
rect -6323 2557 -6277 2603
rect -6203 2557 -6157 2603
rect -6083 2557 -6037 2603
rect -5963 2557 -5917 2603
rect -7163 1597 -7117 1643
rect -7043 1597 -6997 1643
rect -6923 1597 -6877 1643
rect -6803 1597 -6757 1643
rect -6683 1597 -6637 1643
rect -6563 1597 -6517 1643
rect -6443 1597 -6397 1643
rect -6323 1597 -6277 1643
rect -6203 1597 -6157 1643
rect -6083 1597 -6037 1643
rect -5963 1597 -5917 1643
rect -7163 1117 -7117 1163
rect -7043 1117 -6997 1163
rect -6923 1117 -6877 1163
rect -6803 1117 -6757 1163
rect -6683 1117 -6637 1163
rect -6563 1117 -6517 1163
rect -6443 1117 -6397 1163
rect -6323 1117 -6277 1163
rect -6203 1117 -6157 1163
rect -6083 1117 -6037 1163
rect -5963 1117 -5917 1163
rect -7163 637 -7117 683
rect -7043 637 -6997 683
rect -6923 637 -6877 683
rect -6803 637 -6757 683
rect -6683 637 -6637 683
rect -6563 637 -6517 683
rect -6443 637 -6397 683
rect -6323 637 -6277 683
rect -6203 637 -6157 683
rect -6083 637 -6037 683
rect -5963 637 -5917 683
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -6563 -323 -6517 -277
rect -6443 -323 -6397 -277
rect -6323 -323 -6277 -277
rect -6203 -323 -6157 -277
rect -6083 -323 -6037 -277
rect -5963 -323 -5917 -277
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
rect -6563 -1283 -6517 -1237
rect -6443 -1283 -6397 -1237
rect -6323 -1283 -6277 -1237
rect -6203 -1283 -6157 -1237
rect -6083 -1283 -6037 -1237
rect -5963 -1283 -5917 -1237
<< nsubdiffcont >>
rect -7043 3877 -6997 3923
rect -6923 3877 -6877 3923
rect -6803 3877 -6757 3923
rect -6683 3877 -6637 3923
rect -6563 3877 -6517 3923
rect -6443 3877 -6397 3923
rect -6323 3877 -6277 3923
rect -6203 3877 -6157 3923
rect -6083 3877 -6037 3923
rect -7043 2797 -6997 2843
rect -6923 2797 -6877 2843
rect -6803 2797 -6757 2843
rect -6683 2797 -6637 2843
rect -6563 2797 -6517 2843
rect -6443 2797 -6397 2843
rect -6323 2797 -6277 2843
rect -6203 2797 -6157 2843
rect -6083 2797 -6037 2843
<< mvnsubdiffcont >>
rect -7043 5317 -6997 5363
rect -6923 5317 -6877 5363
rect -6803 5317 -6757 5363
rect -6683 5317 -6637 5363
rect -6563 5317 -6517 5363
rect -6443 5317 -6397 5363
rect -6323 5317 -6277 5363
rect -6203 5317 -6157 5363
rect -6083 5317 -6037 5363
rect -7043 4357 -6997 4403
rect -6923 4357 -6877 4403
rect -6803 4357 -6757 4403
rect -6683 4357 -6637 4403
rect -6563 4357 -6517 4403
rect -6443 4357 -6397 4403
rect -6323 4357 -6277 4403
rect -6203 4357 -6157 4403
rect -6083 4357 -6037 4403
<< polysilicon >>
rect -6960 5160 -6840 5220
rect -6720 5160 -6600 5220
rect -6480 5160 -6360 5220
rect -6240 5160 -6120 5220
rect -6960 4680 -6840 4800
rect -6720 4680 -6600 4800
rect -6480 4680 -6360 4800
rect -6240 4680 -6120 4800
rect -6960 4643 -6120 4680
rect -6960 4597 -6923 4643
rect -6877 4597 -6803 4643
rect -6757 4597 -6683 4643
rect -6637 4597 -6563 4643
rect -6517 4597 -6443 4643
rect -6397 4597 -6323 4643
rect -6277 4597 -6203 4643
rect -6157 4597 -6120 4643
rect -6960 4560 -6120 4597
rect -6960 3540 -6840 3600
rect -6720 3540 -6600 3600
rect -6480 3540 -6360 3600
rect -6240 3540 -6120 3600
rect -6960 3120 -6840 3240
rect -6720 3120 -6600 3240
rect -6960 3083 -6600 3120
rect -6960 3037 -6923 3083
rect -6877 3037 -6803 3083
rect -6757 3037 -6683 3083
rect -6637 3037 -6600 3083
rect -6960 3000 -6600 3037
rect -6480 3120 -6360 3240
rect -6240 3120 -6120 3240
rect -6480 3083 -6120 3120
rect -6480 3037 -6443 3083
rect -6397 3037 -6323 3083
rect -6277 3037 -6203 3083
rect -6157 3037 -6120 3083
rect -6480 3000 -6120 3037
rect -6960 -517 -6600 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6803 -517
rect -6757 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -600 -6600 -563
rect -6960 -720 -6840 -600
rect -6720 -720 -6600 -600
rect -6480 -517 -6120 -480
rect -6480 -563 -6443 -517
rect -6397 -563 -6323 -517
rect -6277 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -600 -6120 -563
rect -6480 -720 -6360 -600
rect -6240 -720 -6120 -600
rect -6960 -1140 -6840 -1080
rect -6720 -1140 -6600 -1080
rect -6480 -1140 -6360 -1080
rect -6240 -1140 -6120 -1080
<< polycontact >>
rect -6923 4597 -6877 4643
rect -6803 4597 -6757 4643
rect -6683 4597 -6637 4643
rect -6563 4597 -6517 4643
rect -6443 4597 -6397 4643
rect -6323 4597 -6277 4643
rect -6203 4597 -6157 4643
rect -6923 3037 -6877 3083
rect -6803 3037 -6757 3083
rect -6683 3037 -6637 3083
rect -6443 3037 -6397 3083
rect -6323 3037 -6277 3083
rect -6203 3037 -6157 3083
rect -6923 -563 -6877 -517
rect -6803 -563 -6757 -517
rect -6683 -563 -6637 -517
rect -6443 -563 -6397 -517
rect -6323 -563 -6277 -517
rect -6203 -563 -6157 -517
<< metal1 >>
rect -7200 5603 -5880 5640
rect -7200 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6563 5603
rect -6517 5557 -6443 5603
rect -6397 5557 -6323 5603
rect -6277 5557 -6203 5603
rect -6157 5557 -6083 5603
rect -6037 5557 -5963 5603
rect -5917 5557 -5880 5603
rect -7200 5520 -5880 5557
rect -7200 5366 -5880 5400
rect -7200 5314 -7046 5366
rect -6994 5363 -6566 5366
rect -6514 5363 -6086 5366
rect -6994 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6683 5363
rect -6637 5317 -6566 5363
rect -6514 5317 -6443 5363
rect -6397 5317 -6323 5363
rect -6277 5317 -6203 5363
rect -6157 5317 -6086 5363
rect -6994 5314 -6566 5317
rect -6514 5314 -6086 5317
rect -6034 5314 -5880 5366
rect -7200 5280 -5880 5314
rect -7080 5126 -6960 5160
rect -7080 5074 -7046 5126
rect -6994 5074 -6960 5126
rect -7080 5006 -6960 5074
rect -7080 4954 -7046 5006
rect -6994 4954 -6960 5006
rect -7080 4886 -6960 4954
rect -7080 4834 -7046 4886
rect -6994 4834 -6960 4886
rect -7080 4800 -6960 4834
rect -6840 5126 -6720 5160
rect -6840 5074 -6806 5126
rect -6754 5074 -6720 5126
rect -6840 5006 -6720 5074
rect -6840 4954 -6806 5006
rect -6754 4954 -6720 5006
rect -6840 4886 -6720 4954
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4800 -6720 4834
rect -6600 5126 -6480 5160
rect -6600 5074 -6566 5126
rect -6514 5074 -6480 5126
rect -6600 5006 -6480 5074
rect -6600 4954 -6566 5006
rect -6514 4954 -6480 5006
rect -6600 4886 -6480 4954
rect -6600 4834 -6566 4886
rect -6514 4834 -6480 4886
rect -6600 4800 -6480 4834
rect -6360 5126 -6240 5160
rect -6360 5074 -6326 5126
rect -6274 5074 -6240 5126
rect -6360 5006 -6240 5074
rect -6360 4954 -6326 5006
rect -6274 4954 -6240 5006
rect -6360 4886 -6240 4954
rect -6360 4834 -6326 4886
rect -6274 4834 -6240 4886
rect -6360 4800 -6240 4834
rect -6120 5126 -6000 5160
rect -6120 5074 -6086 5126
rect -6034 5074 -6000 5126
rect -6120 5006 -6000 5074
rect -6120 4954 -6086 5006
rect -6034 4954 -6000 5006
rect -6120 4886 -6000 4954
rect -6120 4834 -6086 4886
rect -6034 4834 -6000 4886
rect -6120 4800 -6000 4834
rect -6960 4646 -6120 4680
rect -6960 4643 -6566 4646
rect -6514 4643 -6120 4646
rect -6960 4597 -6923 4643
rect -6877 4597 -6803 4643
rect -6757 4597 -6683 4643
rect -6637 4597 -6566 4643
rect -6514 4597 -6443 4643
rect -6397 4597 -6323 4643
rect -6277 4597 -6203 4643
rect -6157 4597 -6120 4643
rect -6960 4594 -6566 4597
rect -6514 4594 -6120 4597
rect -6960 4560 -6120 4594
rect -7200 4403 -5880 4440
rect -7200 4357 -7043 4403
rect -6997 4357 -6923 4403
rect -6877 4357 -6803 4403
rect -6757 4357 -6683 4403
rect -6637 4357 -6563 4403
rect -6517 4357 -6443 4403
rect -6397 4357 -6323 4403
rect -6277 4357 -6203 4403
rect -6157 4357 -6083 4403
rect -6037 4357 -5880 4403
rect -7200 4320 -5880 4357
rect -7200 4163 -5880 4200
rect -7200 4117 -7163 4163
rect -7117 4117 -7043 4163
rect -6997 4117 -6923 4163
rect -6877 4117 -6803 4163
rect -6757 4117 -6683 4163
rect -6637 4117 -6563 4163
rect -6517 4117 -6443 4163
rect -6397 4117 -6323 4163
rect -6277 4117 -6203 4163
rect -6157 4117 -6083 4163
rect -6037 4117 -5963 4163
rect -5917 4117 -5880 4163
rect -7200 4080 -5880 4117
rect -7200 3923 -5880 3960
rect -7200 3877 -7043 3923
rect -6997 3877 -6923 3923
rect -6877 3877 -6803 3923
rect -6757 3877 -6683 3923
rect -6637 3877 -6563 3923
rect -6517 3877 -6443 3923
rect -6397 3877 -6323 3923
rect -6277 3877 -6203 3923
rect -6157 3877 -6083 3923
rect -6037 3877 -5880 3923
rect -7200 3840 -5880 3877
rect -7080 3686 -6000 3720
rect -7080 3634 -7046 3686
rect -6994 3634 -6566 3686
rect -6514 3634 -6086 3686
rect -6034 3634 -6000 3686
rect -7080 3600 -6000 3634
rect -7080 3566 -6960 3600
rect -7080 3514 -7046 3566
rect -6994 3514 -6960 3566
rect -6600 3566 -6480 3600
rect -7080 3446 -6960 3514
rect -7080 3394 -7046 3446
rect -6994 3394 -6960 3446
rect -7080 3326 -6960 3394
rect -7080 3274 -7046 3326
rect -6994 3274 -6960 3326
rect -7080 3240 -6960 3274
rect -6840 3446 -6720 3540
rect -6840 3394 -6806 3446
rect -6754 3394 -6720 3446
rect -6840 3326 -6720 3394
rect -6840 3274 -6806 3326
rect -6754 3274 -6720 3326
rect -6840 3240 -6720 3274
rect -6600 3514 -6566 3566
rect -6514 3514 -6480 3566
rect -6120 3566 -6000 3600
rect -6600 3443 -6480 3514
rect -6600 3397 -6563 3443
rect -6517 3397 -6480 3443
rect -6600 3323 -6480 3397
rect -6600 3277 -6563 3323
rect -6517 3277 -6480 3323
rect -6600 3240 -6480 3277
rect -6360 3446 -6240 3540
rect -6360 3394 -6326 3446
rect -6274 3394 -6240 3446
rect -6360 3326 -6240 3394
rect -6360 3274 -6326 3326
rect -6274 3274 -6240 3326
rect -6360 3240 -6240 3274
rect -6120 3514 -6086 3566
rect -6034 3514 -6000 3566
rect -6120 3446 -6000 3514
rect -6120 3394 -6086 3446
rect -6034 3394 -6000 3446
rect -6120 3326 -6000 3394
rect -6120 3274 -6086 3326
rect -6034 3274 -6000 3326
rect -6120 3240 -6000 3274
rect -6960 3086 -6600 3120
rect -6960 3083 -6806 3086
rect -6754 3083 -6600 3086
rect -6960 3037 -6923 3083
rect -6877 3037 -6806 3083
rect -6754 3037 -6683 3083
rect -6637 3037 -6600 3083
rect -6960 3034 -6806 3037
rect -6754 3034 -6600 3037
rect -6960 3000 -6600 3034
rect -6480 3086 -6120 3120
rect -6480 3083 -6326 3086
rect -6274 3083 -6120 3086
rect -6480 3037 -6443 3083
rect -6397 3037 -6326 3083
rect -6274 3037 -6203 3083
rect -6157 3037 -6120 3083
rect -6480 3034 -6326 3037
rect -6274 3034 -6120 3037
rect -6480 3000 -6120 3034
rect -7200 2846 -5880 2880
rect -7200 2794 -7046 2846
rect -6994 2843 -6086 2846
rect -6994 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6683 2843
rect -6637 2797 -6563 2843
rect -6517 2797 -6443 2843
rect -6397 2797 -6323 2843
rect -6277 2797 -6203 2843
rect -6157 2797 -6086 2843
rect -6994 2794 -6086 2797
rect -6034 2794 -5880 2846
rect -7200 2760 -5880 2794
rect -7200 2606 -5880 2640
rect -7200 2603 -7046 2606
rect -6994 2603 -6086 2606
rect -6034 2603 -5880 2606
rect -7200 2557 -7163 2603
rect -7117 2557 -7046 2603
rect -6994 2557 -6923 2603
rect -6877 2557 -6803 2603
rect -6757 2557 -6683 2603
rect -6637 2557 -6563 2603
rect -6517 2557 -6443 2603
rect -6397 2557 -6323 2603
rect -6277 2557 -6203 2603
rect -6157 2557 -6086 2603
rect -6034 2557 -5963 2603
rect -5917 2557 -5880 2603
rect -7200 2554 -7046 2557
rect -6994 2554 -6086 2557
rect -6034 2554 -5880 2557
rect -7200 2520 -5880 2554
rect -7200 1646 -5880 1680
rect -7200 1643 -7046 1646
rect -6994 1643 -6086 1646
rect -6034 1643 -5880 1646
rect -7200 1597 -7163 1643
rect -7117 1597 -7046 1643
rect -6994 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6563 1643
rect -6517 1597 -6443 1643
rect -6397 1597 -6323 1643
rect -6277 1597 -6203 1643
rect -6157 1597 -6086 1643
rect -6034 1597 -5963 1643
rect -5917 1597 -5880 1643
rect -7200 1594 -7046 1597
rect -6994 1594 -6086 1597
rect -6034 1594 -5880 1597
rect -7200 1560 -5880 1594
rect -7200 1166 -5880 1200
rect -7200 1163 -7046 1166
rect -6994 1163 -6086 1166
rect -6034 1163 -5880 1166
rect -7200 1117 -7163 1163
rect -7117 1117 -7046 1163
rect -6994 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6563 1163
rect -6517 1117 -6443 1163
rect -6397 1117 -6323 1163
rect -6277 1117 -6203 1163
rect -6157 1117 -6086 1163
rect -6034 1117 -5963 1163
rect -5917 1117 -5880 1163
rect -7200 1114 -7046 1117
rect -6994 1114 -6086 1117
rect -6034 1114 -5880 1117
rect -7200 1080 -5880 1114
rect -7200 686 -5880 720
rect -7200 683 -7046 686
rect -6994 683 -6086 686
rect -6034 683 -5880 686
rect -7200 637 -7163 683
rect -7117 637 -7046 683
rect -6994 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6563 683
rect -6517 637 -6443 683
rect -6397 637 -6323 683
rect -6277 637 -6203 683
rect -6157 637 -6086 683
rect -6034 637 -5963 683
rect -5917 637 -5880 683
rect -7200 634 -7046 637
rect -6994 634 -6086 637
rect -6034 634 -5880 637
rect -7200 600 -5880 634
rect -7200 -274 -5880 -240
rect -7200 -277 -7046 -274
rect -6994 -277 -6086 -274
rect -6034 -277 -5880 -274
rect -7200 -323 -7163 -277
rect -7117 -323 -7046 -277
rect -6994 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6086 -277
rect -6034 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -326 -7046 -323
rect -6994 -326 -6086 -323
rect -6034 -326 -5880 -323
rect -7200 -360 -5880 -326
rect -6960 -514 -6600 -480
rect -6960 -517 -6806 -514
rect -6754 -517 -6600 -514
rect -6960 -563 -6923 -517
rect -6877 -563 -6806 -517
rect -6754 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -566 -6806 -563
rect -6754 -566 -6600 -563
rect -6960 -600 -6600 -566
rect -6480 -514 -6120 -480
rect -6480 -517 -6326 -514
rect -6274 -517 -6120 -514
rect -6480 -563 -6443 -517
rect -6397 -563 -6326 -517
rect -6274 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -566 -6326 -563
rect -6274 -566 -6120 -563
rect -6480 -600 -6120 -566
rect -7080 -754 -6960 -720
rect -7080 -806 -7046 -754
rect -6994 -806 -6960 -754
rect -7080 -874 -6960 -806
rect -7080 -926 -7046 -874
rect -6994 -926 -6960 -874
rect -7080 -994 -6960 -926
rect -7080 -1046 -7046 -994
rect -6994 -1046 -6960 -994
rect -7080 -1080 -6960 -1046
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -754 -6480 -720
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -754 -6000 -720
rect -6120 -806 -6086 -754
rect -6034 -806 -6000 -754
rect -6120 -874 -6000 -806
rect -6120 -926 -6086 -874
rect -6034 -926 -6000 -874
rect -6120 -994 -6000 -926
rect -6120 -1046 -6086 -994
rect -6034 -1046 -6000 -994
rect -6120 -1080 -6000 -1046
rect -7200 -1234 -5880 -1200
rect -7200 -1237 -7046 -1234
rect -6994 -1237 -6086 -1234
rect -6034 -1237 -5880 -1234
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7046 -1237
rect -6994 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6086 -1237
rect -6034 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1286 -7046 -1283
rect -6994 -1286 -6086 -1283
rect -6034 -1286 -5880 -1283
rect -7200 -1320 -5880 -1286
<< via1 >>
rect -7046 5363 -6994 5366
rect -6566 5363 -6514 5366
rect -6086 5363 -6034 5366
rect -7046 5317 -7043 5363
rect -7043 5317 -6997 5363
rect -6997 5317 -6994 5363
rect -6566 5317 -6563 5363
rect -6563 5317 -6517 5363
rect -6517 5317 -6514 5363
rect -6086 5317 -6083 5363
rect -6083 5317 -6037 5363
rect -6037 5317 -6034 5363
rect -7046 5314 -6994 5317
rect -6566 5314 -6514 5317
rect -6086 5314 -6034 5317
rect -7046 5123 -6994 5126
rect -7046 5077 -7043 5123
rect -7043 5077 -6997 5123
rect -6997 5077 -6994 5123
rect -7046 5074 -6994 5077
rect -7046 5003 -6994 5006
rect -7046 4957 -7043 5003
rect -7043 4957 -6997 5003
rect -6997 4957 -6994 5003
rect -7046 4954 -6994 4957
rect -7046 4883 -6994 4886
rect -7046 4837 -7043 4883
rect -7043 4837 -6997 4883
rect -6997 4837 -6994 4883
rect -7046 4834 -6994 4837
rect -6806 5123 -6754 5126
rect -6806 5077 -6803 5123
rect -6803 5077 -6757 5123
rect -6757 5077 -6754 5123
rect -6806 5074 -6754 5077
rect -6806 5003 -6754 5006
rect -6806 4957 -6803 5003
rect -6803 4957 -6757 5003
rect -6757 4957 -6754 5003
rect -6806 4954 -6754 4957
rect -6806 4883 -6754 4886
rect -6806 4837 -6803 4883
rect -6803 4837 -6757 4883
rect -6757 4837 -6754 4883
rect -6806 4834 -6754 4837
rect -6566 5123 -6514 5126
rect -6566 5077 -6563 5123
rect -6563 5077 -6517 5123
rect -6517 5077 -6514 5123
rect -6566 5074 -6514 5077
rect -6566 5003 -6514 5006
rect -6566 4957 -6563 5003
rect -6563 4957 -6517 5003
rect -6517 4957 -6514 5003
rect -6566 4954 -6514 4957
rect -6566 4883 -6514 4886
rect -6566 4837 -6563 4883
rect -6563 4837 -6517 4883
rect -6517 4837 -6514 4883
rect -6566 4834 -6514 4837
rect -6326 5123 -6274 5126
rect -6326 5077 -6323 5123
rect -6323 5077 -6277 5123
rect -6277 5077 -6274 5123
rect -6326 5074 -6274 5077
rect -6326 5003 -6274 5006
rect -6326 4957 -6323 5003
rect -6323 4957 -6277 5003
rect -6277 4957 -6274 5003
rect -6326 4954 -6274 4957
rect -6326 4883 -6274 4886
rect -6326 4837 -6323 4883
rect -6323 4837 -6277 4883
rect -6277 4837 -6274 4883
rect -6326 4834 -6274 4837
rect -6086 5123 -6034 5126
rect -6086 5077 -6083 5123
rect -6083 5077 -6037 5123
rect -6037 5077 -6034 5123
rect -6086 5074 -6034 5077
rect -6086 5003 -6034 5006
rect -6086 4957 -6083 5003
rect -6083 4957 -6037 5003
rect -6037 4957 -6034 5003
rect -6086 4954 -6034 4957
rect -6086 4883 -6034 4886
rect -6086 4837 -6083 4883
rect -6083 4837 -6037 4883
rect -6037 4837 -6034 4883
rect -6086 4834 -6034 4837
rect -6566 4643 -6514 4646
rect -6566 4597 -6563 4643
rect -6563 4597 -6517 4643
rect -6517 4597 -6514 4643
rect -6566 4594 -6514 4597
rect -7046 3634 -6994 3686
rect -6566 3634 -6514 3686
rect -6086 3634 -6034 3686
rect -7046 3514 -6994 3566
rect -7046 3443 -6994 3446
rect -7046 3397 -7043 3443
rect -7043 3397 -6997 3443
rect -6997 3397 -6994 3443
rect -7046 3394 -6994 3397
rect -7046 3323 -6994 3326
rect -7046 3277 -7043 3323
rect -7043 3277 -6997 3323
rect -6997 3277 -6994 3323
rect -7046 3274 -6994 3277
rect -6806 3443 -6754 3446
rect -6806 3397 -6803 3443
rect -6803 3397 -6757 3443
rect -6757 3397 -6754 3443
rect -6806 3394 -6754 3397
rect -6806 3323 -6754 3326
rect -6806 3277 -6803 3323
rect -6803 3277 -6757 3323
rect -6757 3277 -6754 3323
rect -6806 3274 -6754 3277
rect -6566 3514 -6514 3566
rect -6326 3443 -6274 3446
rect -6326 3397 -6323 3443
rect -6323 3397 -6277 3443
rect -6277 3397 -6274 3443
rect -6326 3394 -6274 3397
rect -6326 3323 -6274 3326
rect -6326 3277 -6323 3323
rect -6323 3277 -6277 3323
rect -6277 3277 -6274 3323
rect -6326 3274 -6274 3277
rect -6086 3514 -6034 3566
rect -6086 3443 -6034 3446
rect -6086 3397 -6083 3443
rect -6083 3397 -6037 3443
rect -6037 3397 -6034 3443
rect -6086 3394 -6034 3397
rect -6086 3323 -6034 3326
rect -6086 3277 -6083 3323
rect -6083 3277 -6037 3323
rect -6037 3277 -6034 3323
rect -6086 3274 -6034 3277
rect -6806 3083 -6754 3086
rect -6806 3037 -6803 3083
rect -6803 3037 -6757 3083
rect -6757 3037 -6754 3083
rect -6806 3034 -6754 3037
rect -6326 3083 -6274 3086
rect -6326 3037 -6323 3083
rect -6323 3037 -6277 3083
rect -6277 3037 -6274 3083
rect -6326 3034 -6274 3037
rect -7046 2843 -6994 2846
rect -6086 2843 -6034 2846
rect -7046 2797 -7043 2843
rect -7043 2797 -6997 2843
rect -6997 2797 -6994 2843
rect -6086 2797 -6083 2843
rect -6083 2797 -6037 2843
rect -6037 2797 -6034 2843
rect -7046 2794 -6994 2797
rect -6086 2794 -6034 2797
rect -7046 2603 -6994 2606
rect -6086 2603 -6034 2606
rect -7046 2557 -7043 2603
rect -7043 2557 -6997 2603
rect -6997 2557 -6994 2603
rect -6086 2557 -6083 2603
rect -6083 2557 -6037 2603
rect -6037 2557 -6034 2603
rect -7046 2554 -6994 2557
rect -6086 2554 -6034 2557
rect -7046 1643 -6994 1646
rect -6086 1643 -6034 1646
rect -7046 1597 -7043 1643
rect -7043 1597 -6997 1643
rect -6997 1597 -6994 1643
rect -6086 1597 -6083 1643
rect -6083 1597 -6037 1643
rect -6037 1597 -6034 1643
rect -7046 1594 -6994 1597
rect -6086 1594 -6034 1597
rect -7046 1163 -6994 1166
rect -6086 1163 -6034 1166
rect -7046 1117 -7043 1163
rect -7043 1117 -6997 1163
rect -6997 1117 -6994 1163
rect -6086 1117 -6083 1163
rect -6083 1117 -6037 1163
rect -6037 1117 -6034 1163
rect -7046 1114 -6994 1117
rect -6086 1114 -6034 1117
rect -7046 683 -6994 686
rect -6086 683 -6034 686
rect -7046 637 -7043 683
rect -7043 637 -6997 683
rect -6997 637 -6994 683
rect -6086 637 -6083 683
rect -6083 637 -6037 683
rect -6037 637 -6034 683
rect -7046 634 -6994 637
rect -6086 634 -6034 637
rect -7046 -277 -6994 -274
rect -6086 -277 -6034 -274
rect -7046 -323 -7043 -277
rect -7043 -323 -6997 -277
rect -6997 -323 -6994 -277
rect -6086 -323 -6083 -277
rect -6083 -323 -6037 -277
rect -6037 -323 -6034 -277
rect -7046 -326 -6994 -323
rect -6086 -326 -6034 -323
rect -6806 -517 -6754 -514
rect -6806 -563 -6803 -517
rect -6803 -563 -6757 -517
rect -6757 -563 -6754 -517
rect -6806 -566 -6754 -563
rect -6326 -517 -6274 -514
rect -6326 -563 -6323 -517
rect -6323 -563 -6277 -517
rect -6277 -563 -6274 -517
rect -6326 -566 -6274 -563
rect -7046 -757 -6994 -754
rect -7046 -803 -7043 -757
rect -7043 -803 -6997 -757
rect -6997 -803 -6994 -757
rect -7046 -806 -6994 -803
rect -7046 -877 -6994 -874
rect -7046 -923 -7043 -877
rect -7043 -923 -6997 -877
rect -6997 -923 -6994 -877
rect -7046 -926 -6994 -923
rect -7046 -997 -6994 -994
rect -7046 -1043 -7043 -997
rect -7043 -1043 -6997 -997
rect -6997 -1043 -6994 -997
rect -7046 -1046 -6994 -1043
rect -6566 -757 -6514 -754
rect -6566 -803 -6563 -757
rect -6563 -803 -6517 -757
rect -6517 -803 -6514 -757
rect -6566 -806 -6514 -803
rect -6566 -877 -6514 -874
rect -6566 -923 -6563 -877
rect -6563 -923 -6517 -877
rect -6517 -923 -6514 -877
rect -6566 -926 -6514 -923
rect -6566 -997 -6514 -994
rect -6566 -1043 -6563 -997
rect -6563 -1043 -6517 -997
rect -6517 -1043 -6514 -997
rect -6566 -1046 -6514 -1043
rect -6086 -757 -6034 -754
rect -6086 -803 -6083 -757
rect -6083 -803 -6037 -757
rect -6037 -803 -6034 -757
rect -6086 -806 -6034 -803
rect -6086 -877 -6034 -874
rect -6086 -923 -6083 -877
rect -6083 -923 -6037 -877
rect -6037 -923 -6034 -877
rect -6086 -926 -6034 -923
rect -6086 -997 -6034 -994
rect -6086 -1043 -6083 -997
rect -6083 -1043 -6037 -997
rect -6037 -1043 -6034 -997
rect -6086 -1046 -6034 -1043
rect -7046 -1237 -6994 -1234
rect -6086 -1237 -6034 -1234
rect -7046 -1283 -7043 -1237
rect -7043 -1283 -6997 -1237
rect -6997 -1283 -6994 -1237
rect -6086 -1283 -6083 -1237
rect -6083 -1283 -6037 -1237
rect -6037 -1283 -6034 -1237
rect -7046 -1286 -6994 -1283
rect -6086 -1286 -6034 -1283
<< metal2 >>
rect -7080 5368 -6960 5400
rect -7080 5312 -7048 5368
rect -6992 5312 -6960 5368
rect -7080 5128 -6960 5312
rect -6600 5368 -6480 5400
rect -6600 5312 -6568 5368
rect -6512 5312 -6480 5368
rect -7080 5072 -7048 5128
rect -6992 5072 -6960 5128
rect -7080 5008 -6960 5072
rect -7080 4952 -7048 5008
rect -6992 4952 -6960 5008
rect -7080 4888 -6960 4952
rect -7080 4832 -7048 4888
rect -6992 4832 -6960 4888
rect -7080 4800 -6960 4832
rect -6840 5126 -6720 5160
rect -6840 5074 -6806 5126
rect -6754 5074 -6720 5126
rect -6840 5006 -6720 5074
rect -6840 4954 -6806 5006
rect -6754 4954 -6720 5006
rect -6840 4886 -6720 4954
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4408 -6720 4834
rect -6600 5128 -6480 5312
rect -6120 5368 -6000 5400
rect -6120 5312 -6088 5368
rect -6032 5312 -6000 5368
rect -6600 5072 -6568 5128
rect -6512 5072 -6480 5128
rect -6600 5008 -6480 5072
rect -6600 4952 -6568 5008
rect -6512 4952 -6480 5008
rect -6600 4888 -6480 4952
rect -6600 4832 -6568 4888
rect -6512 4832 -6480 4888
rect -6600 4800 -6480 4832
rect -6360 5126 -6240 5160
rect -6360 5074 -6326 5126
rect -6274 5074 -6240 5126
rect -6360 5006 -6240 5074
rect -6360 4954 -6326 5006
rect -6274 4954 -6240 5006
rect -6360 4886 -6240 4954
rect -6360 4834 -6326 4886
rect -6274 4834 -6240 4886
rect -6600 4648 -6480 4680
rect -6600 4592 -6568 4648
rect -6512 4592 -6480 4648
rect -6600 4560 -6480 4592
rect -6840 4352 -6808 4408
rect -6752 4352 -6720 4408
rect -7080 3928 -6960 3960
rect -7080 3872 -7048 3928
rect -6992 3872 -6960 3928
rect -7080 3686 -6960 3872
rect -6840 3928 -6720 4352
rect -6360 4408 -6240 4834
rect -6120 5128 -6000 5312
rect -6120 5072 -6088 5128
rect -6032 5072 -6000 5128
rect -6120 5008 -6000 5072
rect -6120 4952 -6088 5008
rect -6032 4952 -6000 5008
rect -6120 4888 -6000 4952
rect -6120 4832 -6088 4888
rect -6032 4832 -6000 4888
rect -6120 4800 -6000 4832
rect -6360 4352 -6328 4408
rect -6272 4352 -6240 4408
rect -6840 3872 -6808 3928
rect -6752 3872 -6720 3928
rect -6840 3840 -6720 3872
rect -6600 3928 -6480 3960
rect -6600 3872 -6568 3928
rect -6512 3872 -6480 3928
rect -7080 3634 -7046 3686
rect -6994 3634 -6960 3686
rect -7080 3566 -6960 3634
rect -7080 3514 -7046 3566
rect -6994 3514 -6960 3566
rect -6600 3686 -6480 3872
rect -6360 3928 -6240 4352
rect -6360 3872 -6328 3928
rect -6272 3872 -6240 3928
rect -6360 3840 -6240 3872
rect -6120 3928 -6000 3960
rect -6120 3872 -6088 3928
rect -6032 3872 -6000 3928
rect -6600 3634 -6566 3686
rect -6514 3634 -6480 3686
rect -6600 3566 -6480 3634
rect -7080 3446 -6960 3514
rect -7080 3394 -7046 3446
rect -6994 3394 -6960 3446
rect -7080 3326 -6960 3394
rect -7080 3274 -7046 3326
rect -6994 3274 -6960 3326
rect -7080 3240 -6960 3274
rect -6840 3446 -6720 3540
rect -6600 3514 -6566 3566
rect -6514 3514 -6480 3566
rect -6120 3686 -6000 3872
rect -6120 3634 -6086 3686
rect -6034 3634 -6000 3686
rect -6120 3566 -6000 3634
rect -6600 3480 -6480 3514
rect -6840 3394 -6806 3446
rect -6754 3394 -6720 3446
rect -6840 3360 -6720 3394
rect -6360 3446 -6240 3540
rect -6360 3394 -6326 3446
rect -6274 3394 -6240 3446
rect -6360 3360 -6240 3394
rect -6840 3326 -6240 3360
rect -6840 3274 -6806 3326
rect -6754 3274 -6326 3326
rect -6274 3274 -6240 3326
rect -6840 3240 -6240 3274
rect -6120 3514 -6086 3566
rect -6034 3514 -6000 3566
rect -6120 3446 -6000 3514
rect -6120 3394 -6086 3446
rect -6034 3394 -6000 3446
rect -6120 3326 -6000 3394
rect -6120 3274 -6086 3326
rect -6034 3274 -6000 3326
rect -6120 3240 -6000 3274
rect -6840 3088 -6720 3120
rect -6840 3032 -6808 3088
rect -6752 3032 -6720 3088
rect -6840 3000 -6720 3032
rect -7080 2848 -6960 2880
rect -7080 2792 -7048 2848
rect -6992 2792 -6960 2848
rect -7080 2760 -6960 2792
rect -7080 2608 -6960 2640
rect -7080 2552 -7048 2608
rect -6992 2552 -6960 2608
rect -7080 1648 -6960 2552
rect -7080 1592 -7048 1648
rect -6992 1592 -6960 1648
rect -7080 1168 -6960 1592
rect -7080 1112 -7048 1168
rect -6992 1112 -6960 1168
rect -7080 688 -6960 1112
rect -7080 632 -7048 688
rect -6992 632 -6960 688
rect -7080 -272 -6960 632
rect -7080 -328 -7048 -272
rect -6992 -328 -6960 -272
rect -7080 -752 -6960 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -7080 -808 -7048 -752
rect -6992 -808 -6960 -752
rect -7080 -872 -6960 -808
rect -7080 -928 -7048 -872
rect -6992 -928 -6960 -872
rect -7080 -992 -6960 -928
rect -7080 -1048 -7048 -992
rect -6992 -1048 -6960 -992
rect -7080 -1232 -6960 -1048
rect -6600 -754 -6480 3240
rect -6360 3088 -6240 3120
rect -6360 3032 -6328 3088
rect -6272 3032 -6240 3088
rect -6360 3000 -6240 3032
rect -6120 2848 -6000 2880
rect -6120 2792 -6088 2848
rect -6032 2792 -6000 2848
rect -6120 2760 -6000 2792
rect -6120 2608 -6000 2640
rect -6120 2552 -6088 2608
rect -6032 2552 -6000 2608
rect -6120 1648 -6000 2552
rect -6120 1592 -6088 1648
rect -6032 1592 -6000 1648
rect -6120 1168 -6000 1592
rect -6120 1112 -6088 1168
rect -6032 1112 -6000 1168
rect -6120 688 -6000 1112
rect -6120 632 -6088 688
rect -6032 632 -6000 688
rect -6120 -272 -6000 632
rect -6120 -328 -6088 -272
rect -6032 -328 -6000 -272
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6120 -752 -6000 -328
rect -6120 -808 -6088 -752
rect -6032 -808 -6000 -752
rect -6120 -872 -6000 -808
rect -6120 -928 -6088 -872
rect -6032 -928 -6000 -872
rect -6120 -992 -6000 -928
rect -6120 -1048 -6088 -992
rect -6032 -1048 -6000 -992
rect -7080 -1288 -7048 -1232
rect -6992 -1288 -6960 -1232
rect -7080 -1320 -6960 -1288
rect -6120 -1232 -6000 -1048
rect -6120 -1288 -6088 -1232
rect -6032 -1288 -6000 -1232
rect -6120 -1320 -6000 -1288
<< via2 >>
rect -7048 5366 -6992 5368
rect -7048 5314 -7046 5366
rect -7046 5314 -6994 5366
rect -6994 5314 -6992 5366
rect -7048 5312 -6992 5314
rect -6568 5366 -6512 5368
rect -6568 5314 -6566 5366
rect -6566 5314 -6514 5366
rect -6514 5314 -6512 5366
rect -6568 5312 -6512 5314
rect -7048 5126 -6992 5128
rect -7048 5074 -7046 5126
rect -7046 5074 -6994 5126
rect -6994 5074 -6992 5126
rect -7048 5072 -6992 5074
rect -7048 5006 -6992 5008
rect -7048 4954 -7046 5006
rect -7046 4954 -6994 5006
rect -6994 4954 -6992 5006
rect -7048 4952 -6992 4954
rect -7048 4886 -6992 4888
rect -7048 4834 -7046 4886
rect -7046 4834 -6994 4886
rect -6994 4834 -6992 4886
rect -7048 4832 -6992 4834
rect -6088 5366 -6032 5368
rect -6088 5314 -6086 5366
rect -6086 5314 -6034 5366
rect -6034 5314 -6032 5366
rect -6088 5312 -6032 5314
rect -6568 5126 -6512 5128
rect -6568 5074 -6566 5126
rect -6566 5074 -6514 5126
rect -6514 5074 -6512 5126
rect -6568 5072 -6512 5074
rect -6568 5006 -6512 5008
rect -6568 4954 -6566 5006
rect -6566 4954 -6514 5006
rect -6514 4954 -6512 5006
rect -6568 4952 -6512 4954
rect -6568 4886 -6512 4888
rect -6568 4834 -6566 4886
rect -6566 4834 -6514 4886
rect -6514 4834 -6512 4886
rect -6568 4832 -6512 4834
rect -6568 4646 -6512 4648
rect -6568 4594 -6566 4646
rect -6566 4594 -6514 4646
rect -6514 4594 -6512 4646
rect -6568 4592 -6512 4594
rect -6808 4352 -6752 4408
rect -7048 3872 -6992 3928
rect -6088 5126 -6032 5128
rect -6088 5074 -6086 5126
rect -6086 5074 -6034 5126
rect -6034 5074 -6032 5126
rect -6088 5072 -6032 5074
rect -6088 5006 -6032 5008
rect -6088 4954 -6086 5006
rect -6086 4954 -6034 5006
rect -6034 4954 -6032 5006
rect -6088 4952 -6032 4954
rect -6088 4886 -6032 4888
rect -6088 4834 -6086 4886
rect -6086 4834 -6034 4886
rect -6034 4834 -6032 4886
rect -6088 4832 -6032 4834
rect -6328 4352 -6272 4408
rect -6808 3872 -6752 3928
rect -6568 3872 -6512 3928
rect -6328 3872 -6272 3928
rect -6088 3872 -6032 3928
rect -6808 3086 -6752 3088
rect -6808 3034 -6806 3086
rect -6806 3034 -6754 3086
rect -6754 3034 -6752 3086
rect -6808 3032 -6752 3034
rect -7048 2846 -6992 2848
rect -7048 2794 -7046 2846
rect -7046 2794 -6994 2846
rect -6994 2794 -6992 2846
rect -7048 2792 -6992 2794
rect -7048 2606 -6992 2608
rect -7048 2554 -7046 2606
rect -7046 2554 -6994 2606
rect -6994 2554 -6992 2606
rect -7048 2552 -6992 2554
rect -7048 1646 -6992 1648
rect -7048 1594 -7046 1646
rect -7046 1594 -6994 1646
rect -6994 1594 -6992 1646
rect -7048 1592 -6992 1594
rect -7048 1166 -6992 1168
rect -7048 1114 -7046 1166
rect -7046 1114 -6994 1166
rect -6994 1114 -6992 1166
rect -7048 1112 -6992 1114
rect -7048 686 -6992 688
rect -7048 634 -7046 686
rect -7046 634 -6994 686
rect -6994 634 -6992 686
rect -7048 632 -6992 634
rect -7048 -274 -6992 -272
rect -7048 -326 -7046 -274
rect -7046 -326 -6994 -274
rect -6994 -326 -6992 -274
rect -7048 -328 -6992 -326
rect -6808 -514 -6752 -512
rect -6808 -566 -6806 -514
rect -6806 -566 -6754 -514
rect -6754 -566 -6752 -514
rect -6808 -568 -6752 -566
rect -7048 -754 -6992 -752
rect -7048 -806 -7046 -754
rect -7046 -806 -6994 -754
rect -6994 -806 -6992 -754
rect -7048 -808 -6992 -806
rect -7048 -874 -6992 -872
rect -7048 -926 -7046 -874
rect -7046 -926 -6994 -874
rect -6994 -926 -6992 -874
rect -7048 -928 -6992 -926
rect -7048 -994 -6992 -992
rect -7048 -1046 -7046 -994
rect -7046 -1046 -6994 -994
rect -6994 -1046 -6992 -994
rect -7048 -1048 -6992 -1046
rect -6328 3086 -6272 3088
rect -6328 3034 -6326 3086
rect -6326 3034 -6274 3086
rect -6274 3034 -6272 3086
rect -6328 3032 -6272 3034
rect -6088 2846 -6032 2848
rect -6088 2794 -6086 2846
rect -6086 2794 -6034 2846
rect -6034 2794 -6032 2846
rect -6088 2792 -6032 2794
rect -6088 2606 -6032 2608
rect -6088 2554 -6086 2606
rect -6086 2554 -6034 2606
rect -6034 2554 -6032 2606
rect -6088 2552 -6032 2554
rect -6088 1646 -6032 1648
rect -6088 1594 -6086 1646
rect -6086 1594 -6034 1646
rect -6034 1594 -6032 1646
rect -6088 1592 -6032 1594
rect -6088 1166 -6032 1168
rect -6088 1114 -6086 1166
rect -6086 1114 -6034 1166
rect -6034 1114 -6032 1166
rect -6088 1112 -6032 1114
rect -6088 686 -6032 688
rect -6088 634 -6086 686
rect -6086 634 -6034 686
rect -6034 634 -6032 686
rect -6088 632 -6032 634
rect -6088 -274 -6032 -272
rect -6088 -326 -6086 -274
rect -6086 -326 -6034 -274
rect -6034 -326 -6032 -274
rect -6088 -328 -6032 -326
rect -6328 -514 -6272 -512
rect -6328 -566 -6326 -514
rect -6326 -566 -6274 -514
rect -6274 -566 -6272 -514
rect -6328 -568 -6272 -566
rect -6088 -754 -6032 -752
rect -6088 -806 -6086 -754
rect -6086 -806 -6034 -754
rect -6034 -806 -6032 -754
rect -6088 -808 -6032 -806
rect -6088 -874 -6032 -872
rect -6088 -926 -6086 -874
rect -6086 -926 -6034 -874
rect -6034 -926 -6032 -874
rect -6088 -928 -6032 -926
rect -6088 -994 -6032 -992
rect -6088 -1046 -6086 -994
rect -6086 -1046 -6034 -994
rect -6034 -1046 -6032 -994
rect -6088 -1048 -6032 -1046
rect -7048 -1234 -6992 -1232
rect -7048 -1286 -7046 -1234
rect -7046 -1286 -6994 -1234
rect -6994 -1286 -6992 -1234
rect -7048 -1288 -6992 -1286
rect -6088 -1234 -6032 -1232
rect -6088 -1286 -6086 -1234
rect -6086 -1286 -6034 -1234
rect -6034 -1286 -6032 -1234
rect -6088 -1288 -6032 -1286
<< metal3 >>
rect -7200 5368 -5880 5400
rect -7200 5312 -7048 5368
rect -6992 5312 -6568 5368
rect -6512 5312 -6088 5368
rect -6032 5312 -5880 5368
rect -7200 5128 -5880 5312
rect -7200 5072 -7048 5128
rect -6992 5072 -6568 5128
rect -6512 5072 -6088 5128
rect -6032 5072 -5880 5128
rect -7200 5008 -5880 5072
rect -7200 4952 -7048 5008
rect -6992 4952 -6568 5008
rect -6512 4952 -6088 5008
rect -6032 4952 -5880 5008
rect -7200 4888 -5880 4952
rect -7200 4832 -7048 4888
rect -6992 4832 -6568 4888
rect -6512 4832 -6088 4888
rect -6032 4832 -5880 4888
rect -7200 4800 -5880 4832
rect -6600 4648 -6480 4680
rect -6600 4592 -6568 4648
rect -6512 4592 -6480 4648
rect -6600 4560 -6480 4592
rect -7200 4408 -5880 4440
rect -7200 4352 -6808 4408
rect -6752 4352 -6328 4408
rect -6272 4352 -5880 4408
rect -7200 4260 -5880 4352
rect -7200 4168 -5880 4200
rect -7200 4112 -6568 4168
rect -6512 4112 -5880 4168
rect -7200 4080 -5880 4112
rect -7200 3928 -5880 4020
rect -7200 3872 -7048 3928
rect -6992 3872 -6808 3928
rect -6752 3872 -6568 3928
rect -6512 3872 -6328 3928
rect -6272 3872 -6088 3928
rect -6032 3872 -5880 3928
rect -7200 3840 -5880 3872
rect -6840 3088 -6720 3120
rect -6840 3032 -6808 3088
rect -6752 3032 -6720 3088
rect -6840 3000 -6720 3032
rect -6360 3088 -6240 3120
rect -6360 3032 -6328 3088
rect -6272 3032 -6240 3088
rect -6360 3000 -6240 3032
rect -7200 2848 -5880 2880
rect -7200 2792 -7048 2848
rect -6992 2792 -6088 2848
rect -6032 2792 -5880 2848
rect -7200 2760 -5880 2792
rect -7200 2608 -5880 2640
rect -7200 2552 -7048 2608
rect -6992 2552 -6088 2608
rect -6032 2552 -5880 2608
rect -7200 2520 -5880 2552
rect -7200 1800 -5880 2400
rect -7200 1648 -5880 1680
rect -7200 1592 -7048 1648
rect -6992 1592 -6088 1648
rect -6032 1592 -5880 1648
rect -7200 1560 -5880 1592
rect -7200 1320 -5880 1440
rect -7200 1168 -5880 1200
rect -7200 1112 -7048 1168
rect -6992 1112 -6088 1168
rect -6032 1112 -5880 1168
rect -7200 1080 -5880 1112
rect -7200 840 -5880 960
rect -7200 688 -5880 720
rect -7200 632 -7048 688
rect -6992 632 -6088 688
rect -6032 632 -5880 688
rect -7200 600 -5880 632
rect -7200 -120 -5880 480
rect -7200 -272 -5880 -240
rect -7200 -328 -7048 -272
rect -6992 -328 -6088 -272
rect -6032 -328 -5880 -272
rect -7200 -360 -5880 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -7200 -752 -5880 -720
rect -7200 -808 -7048 -752
rect -6992 -808 -6088 -752
rect -6032 -808 -5880 -752
rect -7200 -872 -5880 -808
rect -7200 -928 -7048 -872
rect -6992 -928 -6088 -872
rect -6032 -928 -5880 -872
rect -7200 -992 -5880 -928
rect -7200 -1048 -7048 -992
rect -6992 -1048 -6088 -992
rect -6032 -1048 -5880 -992
rect -7200 -1232 -5880 -1048
rect -7200 -1288 -7048 -1232
rect -6992 -1288 -6088 -1232
rect -6032 -1288 -5880 -1232
rect -7200 -1320 -5880 -1288
<< via3 >>
rect -6568 4592 -6512 4648
rect -6808 4352 -6752 4408
rect -6328 4352 -6272 4408
rect -6568 4112 -6512 4168
rect -7048 3872 -6992 3928
rect -6808 3872 -6752 3928
rect -6328 3872 -6272 3928
rect -6088 3872 -6032 3928
rect -6808 3032 -6752 3088
rect -6328 3032 -6272 3088
rect -6808 -568 -6752 -512
rect -6328 -568 -6272 -512
<< metal4 >>
rect -6600 4648 -6480 4680
rect -6600 4592 -6568 4648
rect -6512 4592 -6480 4648
rect -6840 4408 -6720 4440
rect -6840 4352 -6808 4408
rect -6752 4352 -6720 4408
rect -7080 3928 -6960 3960
rect -7080 3872 -7048 3928
rect -6992 3872 -6960 3928
rect -7080 3840 -6960 3872
rect -6840 3928 -6720 4352
rect -6600 4168 -6480 4592
rect -6600 4112 -6568 4168
rect -6512 4112 -6480 4168
rect -6600 4080 -6480 4112
rect -6360 4408 -6240 4440
rect -6360 4352 -6328 4408
rect -6272 4352 -6240 4408
rect -6840 3872 -6808 3928
rect -6752 3872 -6720 3928
rect -6840 3840 -6720 3872
rect -6360 3928 -6240 4352
rect -6360 3872 -6328 3928
rect -6272 3872 -6240 3928
rect -6360 3840 -6240 3872
rect -6120 3928 -6000 3960
rect -6120 3872 -6088 3928
rect -6032 3872 -6000 3928
rect -6120 3840 -6000 3872
rect -6840 3088 -6720 3120
rect -6840 3032 -6808 3088
rect -6752 3032 -6720 3088
rect -6840 2880 -6720 3032
rect -7080 2760 -6720 2880
rect -6840 -512 -6720 2760
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 3088 -6240 3120
rect -6360 3032 -6328 3088
rect -6272 3032 -6240 3088
rect -6360 2880 -6240 3032
rect -6360 2760 -6000 2880
rect -6360 -512 -6240 2760
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
<< labels >>
rlabel metal1 s -6780 -900 -6780 -900 4 dl
rlabel metal1 s -6300 -900 -6300 -900 4 dr
rlabel metal1 s -7020 4140 -7020 4140 4 gnd
rlabel metal1 s -7020 5580 -7020 5580 4 gnd
rlabel metal4 s -6840 -120 -6720 2400 4 inl
port 1 nsew
rlabel metal4 s -6360 -120 -6240 2400 4 inr
port 2 nsew
rlabel metal2 s -6600 -120 -6480 2400 4 out
port 3 nsew
rlabel metal3 s -7200 4800 -5880 5400 4 vdd
port 4 nsew
rlabel metal3 s -7200 4080 -7080 4200 4 gp
port 5 nsew
rlabel metal3 s -7200 2760 -7080 2880 4 bp
port 6 nsew
rlabel metal3 s -7200 4320 -7080 4440 4 vreg
port 7 nsew
rlabel metal3 s -7200 1800 -5880 2400 4 op
port 8 nsew
rlabel metal3 s -7200 1320 -5880 1440 4 im
port 9 nsew
rlabel metal3 s -7200 840 -5880 960 4 ip
port 10 nsew
rlabel metal3 s -7200 -120 -5880 480 4 om
port 11 nsew
rlabel metal3 s -7200 -1320 -5880 -720 4 gnd
port 12 nsew
<< end >>
