magic
tech gf180mcuC
magscale 1 5
timestamp 1665184495
<< metal2 >>
rect -3900 1434 -3840 1440
rect -3900 1146 -3884 1434
rect -3856 1146 -3840 1434
rect -3900 1140 -3840 1146
rect 900 1434 960 1440
rect 900 1146 916 1434
rect 944 1146 960 1434
rect 900 1140 960 1146
rect 1500 1434 1560 1440
rect 1500 1146 1516 1434
rect 1544 1146 1560 1434
rect 1500 1140 1560 1146
rect 6300 1434 6360 1440
rect 6300 1146 6316 1434
rect 6344 1146 6360 1434
rect 6300 1140 6360 1146
rect -2700 704 -2640 720
rect -2700 676 -2684 704
rect -2656 676 -2640 704
rect -2700 660 -2640 676
rect -2100 704 -2040 720
rect -2100 676 -2084 704
rect -2056 676 -2040 704
rect -2100 660 -2040 676
rect 4500 704 4560 720
rect 4500 676 4516 704
rect 4544 676 4560 704
rect 4500 660 4560 676
rect 5100 704 5160 720
rect 5100 676 5116 704
rect 5144 676 5160 704
rect 5100 660 5160 676
rect -1500 464 -1440 480
rect -1500 436 -1484 464
rect -1456 436 -1440 464
rect -1500 420 -1440 436
rect -900 464 -840 480
rect -900 436 -884 464
rect -856 436 -840 464
rect -900 420 -840 436
rect -300 464 -240 480
rect -300 436 -284 464
rect -256 436 -240 464
rect -300 420 -240 436
rect 2700 464 2760 480
rect 2700 436 2716 464
rect 2744 436 2760 464
rect 2700 420 2760 436
rect 3300 464 3360 480
rect 3300 436 3316 464
rect 3344 436 3360 464
rect 3300 420 3360 436
rect 3900 464 3960 480
rect 3900 436 3916 464
rect 3944 436 3960 464
rect 3900 420 3960 436
rect -3300 -6 -3240 0
rect -3300 -294 -3284 -6
rect -3256 -294 -3240 -6
rect -3300 -300 -3240 -294
rect 300 -6 360 0
rect 300 -294 316 -6
rect 344 -294 360 -6
rect 300 -300 360 -294
rect 2100 -6 2160 0
rect 2100 -294 2116 -6
rect 2144 -294 2160 -6
rect 2100 -300 2160 -294
rect 5700 -6 5760 0
rect 5700 -294 5716 -6
rect 5744 -294 5760 -6
rect 5700 -300 5760 -294
<< via2 >>
rect -3884 1146 -3856 1434
rect 916 1146 944 1434
rect 1516 1146 1544 1434
rect 6316 1146 6344 1434
rect -2684 676 -2656 704
rect -2084 676 -2056 704
rect 4516 676 4544 704
rect 5116 676 5144 704
rect -1484 436 -1456 464
rect -884 436 -856 464
rect -284 436 -256 464
rect 2716 436 2744 464
rect 3316 436 3344 464
rect 3916 436 3944 464
rect -3284 -294 -3256 -6
rect 316 -294 344 -6
rect 2116 -294 2144 -6
rect 5716 -294 5744 -6
<< metal3 >>
rect -4680 2640 -4620 2940
rect -4680 2400 -4620 2460
rect -4680 2280 -4620 2340
rect -4680 1620 -4620 1680
rect -4680 1140 -4620 1440
rect -3900 1434 -3840 1440
rect -3900 1146 -3884 1434
rect -3856 1146 -3840 1434
rect -3900 1140 -3840 1146
rect -1980 1434 -1920 1440
rect -1980 1146 -1964 1434
rect -1936 1146 -1920 1434
rect -1980 1140 -1920 1146
rect 900 1434 960 1440
rect 900 1146 916 1434
rect 944 1146 960 1434
rect 900 1140 960 1146
rect 1500 1434 1560 1440
rect 1500 1146 1516 1434
rect 1544 1146 1560 1434
rect 1500 1140 1560 1146
rect 4380 1434 4440 1440
rect 4380 1146 4396 1434
rect 4424 1146 4440 1434
rect 4380 1140 4440 1146
rect 6300 1434 6360 1440
rect 6300 1146 6316 1434
rect 6344 1146 6360 1434
rect 6300 1140 6360 1146
rect -4680 900 -4620 960
rect -4020 944 -3960 960
rect -4020 916 -4004 944
rect -3976 916 -3960 944
rect -4020 900 -3960 916
rect -180 944 -120 960
rect -180 916 -164 944
rect -136 916 -120 944
rect -180 900 -120 916
rect 1020 944 1080 960
rect 1020 916 1036 944
rect 1064 916 1080 944
rect 1020 900 1080 916
rect 1380 944 1440 960
rect 1380 916 1396 944
rect 1424 916 1440 944
rect 1380 900 1440 916
rect 2580 944 2640 960
rect 2580 916 2596 944
rect 2624 916 2640 944
rect 2580 900 2640 916
rect 6420 944 6480 960
rect 6420 916 6436 944
rect 6464 916 6480 944
rect 6420 900 6480 916
rect -4680 660 -4620 720
rect -2700 704 -2640 720
rect -2700 676 -2684 704
rect -2656 676 -2640 704
rect -2700 660 -2640 676
rect -2580 704 -2520 720
rect -2580 676 -2564 704
rect -2536 676 -2520 704
rect -2580 660 -2520 676
rect -2220 704 -2160 720
rect -2220 676 -2204 704
rect -2176 676 -2160 704
rect -2220 660 -2160 676
rect -2100 704 -2040 720
rect -2100 676 -2084 704
rect -2056 676 -2040 704
rect -2100 660 -2040 676
rect -1620 704 -1560 720
rect -1620 676 -1604 704
rect -1576 676 -1560 704
rect -1620 660 -1560 676
rect -780 704 -720 720
rect -780 676 -764 704
rect -736 676 -720 704
rect -780 660 -720 676
rect 3180 704 3240 720
rect 3180 676 3196 704
rect 3224 676 3240 704
rect 3180 660 3240 676
rect 4020 704 4080 720
rect 4020 676 4036 704
rect 4064 676 4080 704
rect 4020 660 4080 676
rect 4500 704 4560 720
rect 4500 676 4516 704
rect 4544 676 4560 704
rect 4500 660 4560 676
rect 4620 704 4680 720
rect 4620 676 4636 704
rect 4664 676 4680 704
rect 4620 660 4680 676
rect 4980 704 5040 720
rect 4980 676 4996 704
rect 5024 676 5040 704
rect 4980 660 5040 676
rect 5100 704 5160 720
rect 5100 676 5116 704
rect 5144 676 5160 704
rect 5100 660 5160 676
rect -4680 420 -4620 480
rect -3780 464 -3720 480
rect -3780 436 -3764 464
rect -3736 436 -3720 464
rect -3780 420 -3720 436
rect -3420 464 -3360 480
rect -3420 436 -3404 464
rect -3376 436 -3360 464
rect -3420 420 -3360 436
rect -1500 464 -1440 480
rect -1500 436 -1484 464
rect -1456 436 -1440 464
rect -1500 420 -1440 436
rect -1380 464 -1320 480
rect -1380 436 -1364 464
rect -1336 436 -1320 464
rect -1380 420 -1320 436
rect -1020 464 -960 480
rect -1020 436 -1004 464
rect -976 436 -960 464
rect -1020 420 -960 436
rect -900 464 -840 480
rect -900 436 -884 464
rect -856 436 -840 464
rect -900 420 -840 436
rect -300 464 -240 480
rect -300 436 -284 464
rect -256 436 -240 464
rect -300 420 -240 436
rect 420 464 480 480
rect 420 436 436 464
rect 464 436 480 464
rect 420 420 480 436
rect 780 464 840 480
rect 780 436 796 464
rect 824 436 840 464
rect 780 420 840 436
rect 1620 464 1680 480
rect 1620 436 1636 464
rect 1664 436 1680 464
rect 1620 420 1680 436
rect 1980 464 2040 480
rect 1980 436 1996 464
rect 2024 436 2040 464
rect 1980 420 2040 436
rect 2700 464 2760 480
rect 2700 436 2716 464
rect 2744 436 2760 464
rect 2700 420 2760 436
rect 3300 464 3360 480
rect 3300 436 3316 464
rect 3344 436 3360 464
rect 3300 420 3360 436
rect 3420 464 3480 480
rect 3420 436 3436 464
rect 3464 436 3480 464
rect 3420 420 3480 436
rect 3780 464 3840 480
rect 3780 436 3796 464
rect 3824 436 3840 464
rect 3780 420 3840 436
rect 3900 464 3960 480
rect 3900 436 3916 464
rect 3944 436 3960 464
rect 3900 420 3960 436
rect 5820 464 5880 480
rect 5820 436 5836 464
rect 5864 436 5880 464
rect 5820 420 5880 436
rect 6180 464 6240 480
rect 6180 436 6196 464
rect 6224 436 6240 464
rect 6180 420 6240 436
rect -4680 180 -4620 240
rect -3180 224 -3120 240
rect -3180 196 -3164 224
rect -3136 196 -3120 224
rect -3180 180 -3120 196
rect -420 224 -360 240
rect -420 196 -404 224
rect -376 196 -360 224
rect -420 180 -360 196
rect 180 224 240 240
rect 180 196 196 224
rect 224 196 240 224
rect 180 180 240 196
rect 2220 224 2280 240
rect 2220 196 2236 224
rect 2264 196 2280 224
rect 2220 180 2280 196
rect 2820 224 2880 240
rect 2820 196 2836 224
rect 2864 196 2880 224
rect 2820 180 2880 196
rect 5580 224 5640 240
rect 5580 196 5596 224
rect 5624 196 5640 224
rect 5580 180 5640 196
rect -4680 -300 -4620 0
rect -3300 -6 -3240 0
rect -3300 -294 -3284 -6
rect -3256 -294 -3240 -6
rect -3300 -300 -3240 -294
rect -2820 -6 -2760 0
rect -2820 -294 -2804 -6
rect -2776 -294 -2760 -6
rect -2820 -300 -2760 -294
rect 300 -6 360 0
rect 300 -294 316 -6
rect 344 -294 360 -6
rect 300 -300 360 -294
rect 2100 -6 2160 0
rect 2100 -294 2116 -6
rect 2144 -294 2160 -6
rect 2100 -300 2160 -294
rect 5220 -6 5280 0
rect 5220 -294 5236 -6
rect 5264 -294 5280 -6
rect 5220 -300 5280 -294
rect 5700 -6 5760 0
rect 5700 -294 5716 -6
rect 5744 -294 5760 -6
rect 5700 -300 5760 -294
rect -4680 -900 -4620 -600
<< via3 >>
rect -1964 1146 -1936 1434
rect 4396 1146 4424 1434
rect -4004 916 -3976 944
rect -164 916 -136 944
rect 1036 916 1064 944
rect 1396 916 1424 944
rect 2596 916 2624 944
rect 6436 916 6464 944
rect -2564 676 -2536 704
rect -2204 676 -2176 704
rect -1604 676 -1576 704
rect -764 676 -736 704
rect 3196 676 3224 704
rect 4036 676 4064 704
rect 4636 676 4664 704
rect 4996 676 5024 704
rect -3764 436 -3736 464
rect -3404 436 -3376 464
rect -1364 436 -1336 464
rect -1004 436 -976 464
rect 436 436 464 464
rect 796 436 824 464
rect 1636 436 1664 464
rect 1996 436 2024 464
rect 3436 436 3464 464
rect 3796 436 3824 464
rect 5836 436 5864 464
rect 6196 436 6224 464
rect -3164 196 -3136 224
rect -404 196 -376 224
rect 196 196 224 224
rect 2236 196 2264 224
rect 2836 196 2864 224
rect 5596 196 5624 224
rect -2804 -294 -2776 -6
rect 5236 -294 5264 -6
<< metal4 >>
rect -1980 1434 -1920 1440
rect -1980 1146 -1964 1434
rect -1936 1146 -1920 1434
rect -1980 1140 -1920 1146
rect 4380 1434 4440 1440
rect 4380 1146 4396 1434
rect 4424 1146 4440 1434
rect 4380 1140 4440 1146
rect -4020 944 -3960 960
rect -4020 916 -4004 944
rect -3976 916 -3960 944
rect -4020 900 -3960 916
rect -180 944 -120 960
rect -180 916 -164 944
rect -136 916 -120 944
rect -180 900 -120 916
rect 1020 944 1080 960
rect 1020 916 1036 944
rect 1064 916 1080 944
rect 1020 900 1080 916
rect 1380 944 1440 960
rect 1380 916 1396 944
rect 1424 916 1440 944
rect 1380 900 1440 916
rect 2580 944 2640 960
rect 2580 916 2596 944
rect 2624 916 2640 944
rect 2580 900 2640 916
rect 6420 944 6480 960
rect 6420 916 6436 944
rect 6464 916 6480 944
rect 6420 900 6480 916
rect -2580 704 -2520 720
rect -2580 676 -2564 704
rect -2536 676 -2520 704
rect -2580 660 -2520 676
rect -2220 704 -2160 720
rect -2220 676 -2204 704
rect -2176 676 -2160 704
rect -2220 660 -2160 676
rect -1620 704 -1560 720
rect -1620 676 -1604 704
rect -1576 676 -1560 704
rect -1620 660 -1560 676
rect -780 704 -720 720
rect -780 676 -764 704
rect -736 676 -720 704
rect -780 660 -720 676
rect 3180 704 3240 720
rect 3180 676 3196 704
rect 3224 676 3240 704
rect 3180 660 3240 676
rect 4020 704 4080 720
rect 4020 676 4036 704
rect 4064 676 4080 704
rect 4020 660 4080 676
rect 4620 704 4680 720
rect 4620 676 4636 704
rect 4664 676 4680 704
rect 4620 660 4680 676
rect 4980 704 5040 720
rect 4980 676 4996 704
rect 5024 676 5040 704
rect 4980 660 5040 676
rect -3780 464 -3720 480
rect -3780 436 -3764 464
rect -3736 436 -3720 464
rect -3780 420 -3720 436
rect -3420 464 -3360 480
rect -3420 436 -3404 464
rect -3376 436 -3360 464
rect -3420 420 -3360 436
rect -1380 464 -1320 480
rect -1380 436 -1364 464
rect -1336 436 -1320 464
rect -1380 420 -1320 436
rect -1020 464 -960 480
rect -1020 436 -1004 464
rect -976 436 -960 464
rect -1020 420 -960 436
rect 420 464 480 480
rect 420 436 436 464
rect 464 436 480 464
rect 420 420 480 436
rect 780 464 840 480
rect 780 436 796 464
rect 824 436 840 464
rect 780 420 840 436
rect 1620 464 1680 480
rect 1620 436 1636 464
rect 1664 436 1680 464
rect 1620 420 1680 436
rect 1980 464 2040 480
rect 1980 436 1996 464
rect 2024 436 2040 464
rect 1980 420 2040 436
rect 3420 464 3480 480
rect 3420 436 3436 464
rect 3464 436 3480 464
rect 3420 420 3480 436
rect 3780 464 3840 480
rect 3780 436 3796 464
rect 3824 436 3840 464
rect 3780 420 3840 436
rect 5820 464 5880 480
rect 5820 436 5836 464
rect 5864 436 5880 464
rect 5820 420 5880 436
rect 6180 464 6240 480
rect 6180 436 6196 464
rect 6224 436 6240 464
rect 6180 420 6240 436
rect -3180 224 -3120 240
rect -3180 196 -3164 224
rect -3136 196 -3120 224
rect -3180 180 -3120 196
rect -420 224 -360 240
rect -420 196 -404 224
rect -376 196 -360 224
rect -420 180 -360 196
rect 180 224 240 240
rect 180 196 196 224
rect 224 196 240 224
rect 180 180 240 196
rect 2220 224 2280 240
rect 2220 196 2236 224
rect 2264 196 2280 224
rect 2220 180 2280 196
rect 2820 224 2880 240
rect 2820 196 2836 224
rect 2864 196 2880 224
rect 2820 180 2880 196
rect 5580 224 5640 240
rect 5580 196 5596 224
rect 5624 196 5640 224
rect 5580 180 5640 196
rect -2820 -6 -2760 0
rect -2820 -294 -2804 -6
rect -2776 -294 -2760 -6
rect -2820 -300 -2760 -294
rect 5220 -6 5280 0
rect 5220 -294 5236 -6
rect 5264 -294 5280 -6
rect 5220 -300 5280 -294
use barthmanf_cell  barthmanf_cell_0
timestamp 1665184495
transform -1 0 3060 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_1
timestamp 1665184495
transform -1 0 2460 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_2
timestamp 1665184495
transform -1 0 1860 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_3
timestamp 1665184495
transform -1 0 1260 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_4
timestamp 1665184495
transform -1 0 660 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_5
timestamp 1665184495
transform -1 0 60 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_6
timestamp 1665184495
transform -1 0 -540 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_7
timestamp 1665184495
transform -1 0 -1140 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_8
timestamp 1665184495
transform -1 0 -1740 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_9
timestamp 1665184495
transform 1 0 4200 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_10
timestamp 1665184495
transform 1 0 3600 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_11
timestamp 1665184495
transform 1 0 3000 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_12
timestamp 1665184495
transform 1 0 2400 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_13
timestamp 1665184495
transform 1 0 1800 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_14
timestamp 1665184495
transform 1 0 1200 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_15
timestamp 1665184495
transform 1 0 600 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_16
timestamp 1665184495
transform 1 0 0 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_cell  barthmanf_cell_17
timestamp 1665184495
transform 1 0 -600 0 1 -240
box -3600 -660 -2940 3300
use barthmanf_edge  barthmanf_edge_0
timestamp 1665184495
transform -1 0 3300 0 1 -240
box -3780 -660 -3300 3300
use barthmanf_edge  barthmanf_edge_1
timestamp 1665184495
transform 1 0 -840 0 1 -240
box -3780 -660 -3300 3300
<< labels >>
rlabel metal3 s -4650 690 -4650 690 4 x
rlabel metal3 s -4650 450 -4650 450 4 y
rlabel metal3 s -4680 180 -4620 240 4 ip
port 1 nsew
rlabel metal3 s -4680 900 -4620 960 4 im
port 2 nsew
rlabel metal3 s -4680 1140 -4620 1440 4 op
port 3 nsew
rlabel metal3 s -4680 -300 -4620 0 4 om
port 4 nsew
rlabel metal3 s -4680 2640 -4620 2940 4 vdd
port 5 nsew
rlabel metal3 s -4680 2280 -4620 2340 4 gp
port 6 nsew
rlabel metal3 s -4680 1620 -4620 1680 4 bp
port 7 nsew
rlabel metal3 s -4680 2400 -4620 2460 4 vreg
port 8 nsew
rlabel metal3 s -4680 -900 -4620 -600 4 gnd
port 9 nsew
<< end >>
