magic
tech gf180mcuC
magscale 1 5
timestamp 1665299795
<< error_s >>
rect -5062 3962 -4598 3982
rect -5062 3954 -5042 3962
rect -5034 3954 -5006 3962
rect -4958 3954 -4930 3962
rect -4882 3954 -4854 3962
rect -4806 3954 -4778 3962
rect -4730 3954 -4702 3962
rect -4654 3954 -4626 3962
rect -4618 3954 -4598 3962
rect -5034 3926 -4986 3954
rect -4958 3926 -4910 3954
rect -4882 3926 -4834 3954
rect -4806 3926 -4758 3954
rect -4730 3926 -4682 3954
rect -4654 3926 -4598 3954
rect -5062 3878 -5042 3906
rect -5034 3878 -5006 3898
rect -4958 3878 -4930 3898
rect -4882 3878 -4854 3898
rect -4806 3878 -4778 3898
rect -4730 3878 -4702 3898
rect -4654 3878 -4626 3898
rect -4618 3878 -4598 3906
rect -5034 3850 -4986 3878
rect -4958 3850 -4910 3878
rect -4882 3850 -4834 3878
rect -4806 3850 -4758 3878
rect -4730 3850 -4682 3878
rect -4654 3850 -4598 3878
rect -5062 3802 -5042 3830
rect -5034 3802 -5006 3822
rect -4958 3802 -4930 3822
rect -4882 3802 -4854 3822
rect -4806 3802 -4778 3822
rect -4730 3802 -4702 3822
rect -4654 3802 -4626 3822
rect -4618 3802 -4598 3830
rect -5034 3774 -4986 3802
rect -4958 3774 -4910 3802
rect -4882 3774 -4834 3802
rect -4806 3774 -4758 3802
rect -4730 3774 -4682 3802
rect -4654 3774 -4598 3802
rect -5062 3726 -5042 3754
rect -5034 3726 -5006 3746
rect -4958 3726 -4930 3746
rect -4882 3726 -4854 3746
rect -4806 3726 -4778 3746
rect -4730 3726 -4702 3746
rect -4654 3726 -4626 3746
rect -4618 3726 -4598 3754
rect -5034 3698 -4986 3726
rect -4958 3698 -4910 3726
rect -4882 3698 -4834 3726
rect -4806 3698 -4758 3726
rect -4730 3698 -4682 3726
rect -4654 3698 -4598 3726
rect -5062 3650 -5042 3678
rect -5034 3650 -5006 3670
rect -4958 3650 -4930 3670
rect -4882 3650 -4854 3670
rect -4806 3650 -4778 3670
rect -4730 3650 -4702 3670
rect -4654 3650 -4626 3670
rect -4618 3650 -4598 3678
rect -5034 3622 -4986 3650
rect -4958 3622 -4910 3650
rect -4882 3622 -4834 3650
rect -4806 3622 -4758 3650
rect -4730 3622 -4682 3650
rect -4654 3622 -4598 3650
rect -5062 3574 -5042 3602
rect -5034 3574 -5006 3594
rect -4958 3574 -4930 3594
rect -4882 3574 -4854 3594
rect -4806 3574 -4778 3594
rect -4730 3574 -4702 3594
rect -4654 3574 -4626 3594
rect -4618 3574 -4598 3602
rect -5034 3546 -4986 3574
rect -4958 3546 -4910 3574
rect -4882 3546 -4834 3574
rect -4806 3546 -4758 3574
rect -4730 3546 -4682 3574
rect -4654 3546 -4598 3574
rect -5062 -1258 -4598 -1238
rect -5062 -1266 -5042 -1258
rect -5034 -1266 -5006 -1258
rect -4958 -1266 -4930 -1258
rect -4882 -1266 -4854 -1258
rect -4806 -1266 -4778 -1258
rect -4730 -1266 -4702 -1258
rect -4654 -1266 -4626 -1258
rect -4618 -1266 -4598 -1258
rect -5034 -1294 -4986 -1266
rect -4958 -1294 -4910 -1266
rect -4882 -1294 -4834 -1266
rect -4806 -1294 -4758 -1266
rect -4730 -1294 -4682 -1266
rect -4654 -1294 -4598 -1266
rect -5062 -1342 -5042 -1314
rect -5034 -1342 -5006 -1322
rect -4958 -1342 -4930 -1322
rect -4882 -1342 -4854 -1322
rect -4806 -1342 -4778 -1322
rect -4730 -1342 -4702 -1322
rect -4654 -1342 -4626 -1322
rect -4618 -1342 -4598 -1314
rect -5034 -1370 -4986 -1342
rect -4958 -1370 -4910 -1342
rect -4882 -1370 -4834 -1342
rect -4806 -1370 -4758 -1342
rect -4730 -1370 -4682 -1342
rect -4654 -1370 -4598 -1342
rect -5062 -1418 -5042 -1390
rect -5034 -1418 -5006 -1398
rect -4958 -1418 -4930 -1398
rect -4882 -1418 -4854 -1398
rect -4806 -1418 -4778 -1398
rect -4730 -1418 -4702 -1398
rect -4654 -1418 -4626 -1398
rect -4618 -1418 -4598 -1390
rect -5034 -1446 -4986 -1418
rect -4958 -1446 -4910 -1418
rect -4882 -1446 -4834 -1418
rect -4806 -1446 -4758 -1418
rect -4730 -1446 -4682 -1418
rect -4654 -1446 -4598 -1418
rect -5062 -1494 -5042 -1466
rect -5034 -1494 -5006 -1474
rect -4958 -1494 -4930 -1474
rect -4882 -1494 -4854 -1474
rect -4806 -1494 -4778 -1474
rect -4730 -1494 -4702 -1474
rect -4654 -1494 -4626 -1474
rect -4618 -1494 -4598 -1466
rect -5034 -1522 -4986 -1494
rect -4958 -1522 -4910 -1494
rect -4882 -1522 -4834 -1494
rect -4806 -1522 -4758 -1494
rect -4730 -1522 -4682 -1494
rect -4654 -1522 -4598 -1494
rect -5062 -1570 -5042 -1542
rect -5034 -1570 -5006 -1550
rect -4958 -1570 -4930 -1550
rect -4882 -1570 -4854 -1550
rect -4806 -1570 -4778 -1550
rect -4730 -1570 -4702 -1550
rect -4654 -1570 -4626 -1550
rect -4618 -1570 -4598 -1542
rect -5034 -1598 -4986 -1570
rect -4958 -1598 -4910 -1570
rect -4882 -1598 -4834 -1570
rect -4806 -1598 -4758 -1570
rect -4730 -1598 -4682 -1570
rect -4654 -1598 -4598 -1570
rect -5062 -1646 -5042 -1618
rect -5034 -1646 -5006 -1626
rect -4958 -1646 -4930 -1626
rect -4882 -1646 -4854 -1626
rect -4806 -1646 -4778 -1626
rect -4730 -1646 -4702 -1626
rect -4654 -1646 -4626 -1626
rect -4618 -1646 -4598 -1618
rect -5034 -1674 -4986 -1646
rect -4958 -1674 -4910 -1646
rect -4882 -1674 -4834 -1646
rect -4806 -1674 -4758 -1646
rect -4730 -1674 -4682 -1646
rect -4654 -1674 -4598 -1646
<< metal2 >>
rect -1440 1480 -1380 1500
rect -1440 1400 -1424 1480
rect -1396 1400 -1380 1480
rect -1440 1380 -1380 1400
rect 1560 1480 1620 1500
rect 1560 1400 1576 1480
rect 1604 1400 1620 1480
rect 1560 1380 1620 1400
rect 3360 1480 3420 1500
rect 3360 1400 3376 1480
rect 3404 1400 3420 1480
rect 3360 1380 3420 1400
rect 3960 1480 4020 1500
rect 3960 1400 3976 1480
rect 4004 1400 4020 1480
rect 3960 1380 4020 1400
rect 5760 1480 5820 1500
rect 5760 1400 5776 1480
rect 5804 1400 5820 1480
rect 5760 1380 5820 1400
rect 6360 1480 6420 1500
rect 6360 1400 6376 1480
rect 6404 1400 6420 1480
rect 6360 1380 6420 1400
rect 8160 1480 8220 1500
rect 8160 1400 8176 1480
rect 8204 1400 8220 1480
rect 8160 1380 8220 1400
rect 11160 1480 11220 1500
rect 11160 1400 11176 1480
rect 11204 1400 11220 1480
rect 11160 1380 11220 1400
rect -4440 1304 -4380 1320
rect -4440 1276 -4424 1304
rect -4396 1276 -4380 1304
rect -4440 1260 -4380 1276
rect -3840 1304 -3780 1320
rect -3840 1276 -3824 1304
rect -3796 1276 -3780 1304
rect -3840 1260 -3780 1276
rect 960 1304 1020 1320
rect 960 1276 976 1304
rect 1004 1276 1020 1304
rect 960 1260 1020 1276
rect 8760 1304 8820 1320
rect 8760 1276 8776 1304
rect 8804 1276 8820 1304
rect 8760 1260 8820 1276
rect 13560 1304 13620 1320
rect 13560 1276 13576 1304
rect 13604 1276 13620 1304
rect 13560 1260 13620 1276
rect 14160 1304 14220 1320
rect 14160 1276 14176 1304
rect 14204 1276 14220 1304
rect 14160 1260 14220 1276
rect -1440 1180 -1380 1200
rect -1440 1100 -1424 1180
rect -1396 1100 -1380 1180
rect -1440 1080 -1380 1100
rect 1560 1180 1620 1200
rect 1560 1100 1576 1180
rect 1604 1100 1620 1180
rect 1560 1080 1620 1100
rect 3360 1180 3420 1200
rect 3360 1100 3376 1180
rect 3404 1100 3420 1180
rect 3360 1080 3420 1100
rect 3960 1180 4020 1200
rect 3960 1100 3976 1180
rect 4004 1100 4020 1180
rect 3960 1080 4020 1100
rect 5760 1180 5820 1200
rect 5760 1100 5776 1180
rect 5804 1100 5820 1180
rect 5760 1080 5820 1100
rect 6360 1180 6420 1200
rect 6360 1100 6376 1180
rect 6404 1100 6420 1180
rect 6360 1080 6420 1100
rect 8160 1180 8220 1200
rect 8160 1100 8176 1180
rect 8204 1100 8220 1180
rect 8160 1080 8220 1100
rect 11160 1180 11220 1200
rect 11160 1100 11176 1180
rect 11204 1100 11220 1180
rect 11160 1080 11220 1100
rect -840 644 -780 660
rect -840 616 -824 644
rect -796 616 -780 644
rect -840 600 -780 616
rect -240 644 -180 660
rect -240 616 -224 644
rect -196 616 -180 644
rect -240 600 -180 616
rect 9960 644 10020 660
rect 9960 616 9976 644
rect 10004 616 10020 644
rect 9960 600 10020 616
rect 10560 644 10620 660
rect 10560 616 10576 644
rect 10604 616 10620 644
rect 10560 600 10620 616
rect -2040 160 -1980 180
rect -2040 80 -2024 160
rect -1996 80 -1980 160
rect -2040 60 -1980 80
rect 2160 160 2220 180
rect 2160 80 2176 160
rect 2204 80 2220 160
rect 2160 60 2220 80
rect 2760 160 2820 180
rect 2760 80 2776 160
rect 2804 80 2820 160
rect 2760 60 2820 80
rect 4560 160 4620 180
rect 4560 80 4576 160
rect 4604 80 4620 160
rect 4560 60 4620 80
rect 5160 160 5220 180
rect 5160 80 5176 160
rect 5204 80 5220 160
rect 5160 60 5220 80
rect 6960 160 7020 180
rect 6960 80 6976 160
rect 7004 80 7020 160
rect 6960 60 7020 80
rect 7560 160 7620 180
rect 7560 80 7576 160
rect 7604 80 7620 160
rect 7560 60 7620 80
rect 11760 160 11820 180
rect 11760 80 11776 160
rect 11804 80 11820 160
rect 11760 60 11820 80
rect -3240 -16 -3180 0
rect -3240 -44 -3224 -16
rect -3196 -44 -3180 -16
rect -3240 -60 -3180 -44
rect -2640 -16 -2580 0
rect -2640 -44 -2624 -16
rect -2596 -44 -2580 -16
rect -2640 -60 -2580 -44
rect 360 -16 420 0
rect 360 -44 376 -16
rect 404 -44 420 -16
rect 360 -60 420 -44
rect 9360 -16 9420 0
rect 9360 -44 9376 -16
rect 9404 -44 9420 -16
rect 9360 -60 9420 -44
rect 12360 -16 12420 0
rect 12360 -44 12376 -16
rect 12404 -44 12420 -16
rect 12360 -60 12420 -44
rect 12960 -16 13020 0
rect 12960 -44 12976 -16
rect 13004 -44 13020 -16
rect 12960 -60 13020 -44
rect -2040 -140 -1980 -120
rect -2040 -220 -2024 -140
rect -1996 -220 -1980 -140
rect -2040 -240 -1980 -220
rect 2160 -140 2220 -120
rect 2160 -220 2176 -140
rect 2204 -220 2220 -140
rect 2160 -240 2220 -220
rect 2760 -140 2820 -120
rect 2760 -220 2776 -140
rect 2804 -220 2820 -140
rect 2760 -240 2820 -220
rect 4560 -140 4620 -120
rect 4560 -220 4576 -140
rect 4604 -220 4620 -140
rect 4560 -240 4620 -220
rect 5160 -140 5220 -120
rect 5160 -220 5176 -140
rect 5204 -220 5220 -140
rect 5160 -240 5220 -220
rect 6960 -140 7020 -120
rect 6960 -220 6976 -140
rect 7004 -220 7020 -140
rect 6960 -240 7020 -220
rect 7560 -140 7620 -120
rect 7560 -220 7576 -140
rect 7604 -220 7620 -140
rect 7560 -240 7620 -220
rect 11760 -140 11820 -120
rect 11760 -220 11776 -140
rect 11804 -220 11820 -140
rect 11760 -240 11820 -220
<< via2 >>
rect -1424 1400 -1396 1480
rect 1576 1400 1604 1480
rect 3376 1400 3404 1480
rect 3976 1400 4004 1480
rect 5776 1400 5804 1480
rect 6376 1400 6404 1480
rect 8176 1400 8204 1480
rect 11176 1400 11204 1480
rect -4424 1276 -4396 1304
rect -3824 1276 -3796 1304
rect 976 1276 1004 1304
rect 8776 1276 8804 1304
rect 13576 1276 13604 1304
rect 14176 1276 14204 1304
rect -1424 1100 -1396 1180
rect 1576 1100 1604 1180
rect 3376 1100 3404 1180
rect 3976 1100 4004 1180
rect 5776 1100 5804 1180
rect 6376 1100 6404 1180
rect 8176 1100 8204 1180
rect 11176 1100 11204 1180
rect -824 616 -796 644
rect -224 616 -196 644
rect 9976 616 10004 644
rect 10576 616 10604 644
rect -2024 80 -1996 160
rect 2176 80 2204 160
rect 2776 80 2804 160
rect 4576 80 4604 160
rect 5176 80 5204 160
rect 6976 80 7004 160
rect 7576 80 7604 160
rect 11776 80 11804 160
rect -3224 -44 -3196 -16
rect -2624 -44 -2596 -16
rect 376 -44 404 -16
rect 9376 -44 9404 -16
rect 12376 -44 12404 -16
rect 12976 -44 13004 -16
rect -2024 -220 -1996 -140
rect 2176 -220 2204 -140
rect 2776 -220 2804 -140
rect 4576 -220 4604 -140
rect 5176 -220 5204 -140
rect 6976 -220 7004 -140
rect 7576 -220 7604 -140
rect 11776 -220 11804 -140
<< mimcap >>
rect -5100 3962 14880 4200
rect -5100 3538 -5042 3962
rect -4618 3538 14880 3962
rect -5100 3480 14880 3538
rect -5100 -1258 14880 -1200
rect -5100 -1682 -5042 -1258
rect -4618 -1682 14880 -1258
rect -5100 -1920 14880 -1682
<< mimcapcontact >>
rect -5042 3538 -4618 3962
rect -5042 -1682 -4618 -1258
<< metal3 >>
rect -5220 2700 -5160 3000
rect -5220 2430 -5160 2520
rect -5220 2340 -5160 2400
rect -5220 1680 -5160 1740
rect -5520 1465 -5160 1500
rect -5520 1385 -5504 1465
rect -5476 1385 -5264 1465
rect -5236 1385 -5160 1465
rect -5520 1350 -5160 1385
rect -1440 1480 -1380 1500
rect -1440 1400 -1424 1480
rect -1396 1400 -1380 1480
rect -1440 1380 -1380 1400
rect -120 1480 -60 1500
rect -120 1400 -104 1480
rect -76 1400 -60 1480
rect -120 1380 -60 1400
rect 1560 1480 1620 1500
rect 1560 1400 1576 1480
rect 1604 1400 1620 1480
rect 1560 1380 1620 1400
rect 3360 1480 3420 1500
rect 3360 1400 3376 1480
rect 3404 1400 3420 1480
rect 3360 1380 3420 1400
rect 3960 1480 4020 1500
rect 3960 1400 3976 1480
rect 4004 1400 4020 1480
rect 3960 1380 4020 1400
rect 5760 1480 5820 1500
rect 5760 1400 5776 1480
rect 5804 1400 5820 1480
rect 5760 1380 5820 1400
rect 6360 1480 6420 1500
rect 6360 1400 6376 1480
rect 6404 1400 6420 1480
rect 6360 1380 6420 1400
rect 8160 1480 8220 1500
rect 8160 1400 8176 1480
rect 8204 1400 8220 1480
rect 8160 1380 8220 1400
rect 9840 1480 9900 1500
rect 9840 1400 9856 1480
rect 9884 1400 9900 1480
rect 9840 1380 9900 1400
rect 11160 1480 11220 1500
rect 11160 1400 11176 1480
rect 11204 1400 11220 1480
rect 11160 1380 11220 1400
rect -5520 1304 -5160 1320
rect -5520 1276 -5384 1304
rect -5356 1276 -5160 1304
rect -5520 1260 -5160 1276
rect -4440 1304 -4380 1320
rect -4440 1276 -4424 1304
rect -4396 1276 -4380 1304
rect -4440 1260 -4380 1276
rect -4320 1304 -4260 1320
rect -4320 1276 -4304 1304
rect -4276 1276 -4260 1304
rect -4320 1260 -4260 1276
rect -3840 1304 -3780 1320
rect -3840 1276 -3824 1304
rect -3796 1276 -3780 1304
rect -3840 1260 -3780 1276
rect -3360 1304 -3300 1320
rect -3360 1276 -3344 1304
rect -3316 1276 -3300 1304
rect -3360 1260 -3300 1276
rect -1560 1304 -1500 1320
rect -1560 1276 -1544 1304
rect -1516 1276 -1500 1304
rect -1560 1260 -1500 1276
rect -1320 1304 -1260 1320
rect -1320 1276 -1304 1304
rect -1276 1276 -1260 1304
rect -1320 1260 -1260 1276
rect 960 1304 1020 1320
rect 960 1276 976 1304
rect 1004 1276 1020 1304
rect 960 1260 1020 1276
rect 1440 1304 1500 1320
rect 1440 1276 1456 1304
rect 1484 1276 1500 1304
rect 1440 1260 1500 1276
rect 1680 1304 1740 1320
rect 1680 1276 1696 1304
rect 1724 1276 1740 1304
rect 1680 1260 1740 1276
rect 8040 1304 8100 1320
rect 8040 1276 8056 1304
rect 8084 1276 8100 1304
rect 8040 1260 8100 1276
rect 8280 1304 8340 1320
rect 8280 1276 8296 1304
rect 8324 1276 8340 1304
rect 8280 1260 8340 1276
rect 8760 1304 8820 1320
rect 8760 1276 8776 1304
rect 8804 1276 8820 1304
rect 8760 1260 8820 1276
rect 11040 1304 11100 1320
rect 11040 1276 11056 1304
rect 11084 1276 11100 1304
rect 11040 1260 11100 1276
rect 11280 1304 11340 1320
rect 11280 1276 11296 1304
rect 11324 1276 11340 1304
rect 11280 1260 11340 1276
rect 13080 1304 13140 1320
rect 13080 1276 13096 1304
rect 13124 1276 13140 1304
rect 13080 1260 13140 1276
rect 13560 1304 13620 1320
rect 13560 1276 13576 1304
rect 13604 1276 13620 1304
rect 13560 1260 13620 1276
rect 14040 1304 14100 1320
rect 14040 1276 14056 1304
rect 14084 1276 14100 1304
rect 14040 1260 14100 1276
rect 14160 1304 14220 1320
rect 14160 1276 14176 1304
rect 14204 1276 14220 1304
rect 14160 1260 14220 1276
rect -5520 1195 -5160 1230
rect -5520 1115 -5504 1195
rect -5476 1115 -5264 1195
rect -5236 1115 -5160 1195
rect -5520 1080 -5160 1115
rect -1440 1180 -1380 1200
rect -1440 1100 -1424 1180
rect -1396 1100 -1380 1180
rect -1440 1080 -1380 1100
rect -120 1180 -60 1200
rect -120 1100 -104 1180
rect -76 1100 -60 1180
rect -120 1080 -60 1100
rect 1560 1180 1620 1200
rect 1560 1100 1576 1180
rect 1604 1100 1620 1180
rect 1560 1080 1620 1100
rect 3360 1180 3420 1200
rect 3360 1100 3376 1180
rect 3404 1100 3420 1180
rect 3360 1080 3420 1100
rect 3960 1180 4020 1200
rect 3960 1100 3976 1180
rect 4004 1100 4020 1180
rect 3960 1080 4020 1100
rect 5760 1180 5820 1200
rect 5760 1100 5776 1180
rect 5804 1100 5820 1180
rect 5760 1080 5820 1100
rect 6360 1180 6420 1200
rect 6360 1100 6376 1180
rect 6404 1100 6420 1180
rect 6360 1080 6420 1100
rect 8160 1180 8220 1200
rect 8160 1100 8176 1180
rect 8204 1100 8220 1180
rect 8160 1080 8220 1100
rect 9840 1180 9900 1200
rect 9840 1100 9856 1180
rect 9884 1100 9900 1180
rect 9840 1080 9900 1100
rect 11160 1180 11220 1200
rect 11160 1100 11176 1180
rect 11204 1100 11220 1180
rect 11160 1080 11220 1100
rect -5220 840 -5160 900
rect -3120 884 -3060 900
rect -3120 856 -3104 884
rect -3076 856 -3060 884
rect -3120 840 -3060 856
rect -2520 884 -2460 900
rect -2520 856 -2504 884
rect -2476 856 -2460 884
rect -2520 840 -2460 856
rect 3240 884 3300 900
rect 3240 856 3256 884
rect 3284 856 3300 884
rect 3240 840 3300 856
rect 3480 884 3540 900
rect 3480 856 3496 884
rect 3524 856 3540 884
rect 3480 840 3540 856
rect 3840 884 3900 900
rect 3840 856 3856 884
rect 3884 856 3900 884
rect 3840 840 3900 856
rect 4080 884 4140 900
rect 4080 856 4096 884
rect 4124 856 4140 884
rect 4080 840 4140 856
rect 5640 884 5700 900
rect 5640 856 5656 884
rect 5684 856 5700 884
rect 5640 840 5700 856
rect 5880 884 5940 900
rect 5880 856 5896 884
rect 5924 856 5940 884
rect 5880 840 5940 856
rect 6240 884 6300 900
rect 6240 856 6256 884
rect 6284 856 6300 884
rect 6240 840 6300 856
rect 6480 884 6540 900
rect 6480 856 6496 884
rect 6524 856 6540 884
rect 6480 840 6540 856
rect 12240 884 12300 900
rect 12240 856 12256 884
rect 12284 856 12300 884
rect 12240 840 12300 856
rect 12840 884 12900 900
rect 12840 856 12856 884
rect 12884 856 12900 884
rect 12840 840 12900 856
rect -5220 600 -5160 660
rect -840 644 -780 660
rect -840 616 -824 644
rect -796 616 -780 644
rect -840 600 -780 616
rect -720 644 -660 660
rect -720 616 -704 644
rect -676 616 -660 644
rect -720 600 -660 616
rect -360 644 -300 660
rect -360 616 -344 644
rect -316 616 -300 644
rect -360 600 -300 616
rect -240 644 -180 660
rect -240 616 -224 644
rect -196 616 -180 644
rect -240 600 -180 616
rect 240 644 300 660
rect 240 616 256 644
rect 284 616 300 644
rect 240 600 300 616
rect 480 644 540 660
rect 480 616 496 644
rect 524 616 540 644
rect 480 600 540 616
rect 840 644 900 660
rect 840 616 856 644
rect 884 616 900 644
rect 840 600 900 616
rect 1080 644 1140 660
rect 1080 616 1096 644
rect 1124 616 1140 644
rect 1080 600 1140 616
rect 8640 644 8700 660
rect 8640 616 8656 644
rect 8684 616 8700 644
rect 8640 600 8700 616
rect 8880 644 8940 660
rect 8880 616 8896 644
rect 8924 616 8940 644
rect 8880 600 8940 616
rect 9240 644 9300 660
rect 9240 616 9256 644
rect 9284 616 9300 644
rect 9240 600 9300 616
rect 9480 644 9540 660
rect 9480 616 9496 644
rect 9524 616 9540 644
rect 9480 600 9540 616
rect 9960 644 10020 660
rect 9960 616 9976 644
rect 10004 616 10020 644
rect 9960 600 10020 616
rect 10080 644 10140 660
rect 10080 616 10096 644
rect 10124 616 10140 644
rect 10080 600 10140 616
rect 10440 644 10500 660
rect 10440 616 10456 644
rect 10484 616 10500 644
rect 10440 600 10500 616
rect 10560 644 10620 660
rect 10560 616 10576 644
rect 10604 616 10620 644
rect 10560 600 10620 616
rect -5220 360 -5160 420
rect -4560 404 -4500 420
rect -4560 376 -4544 404
rect -4516 376 -4500 404
rect -4560 360 -4500 376
rect -3960 404 -3900 420
rect -3960 376 -3944 404
rect -3916 376 -3900 404
rect -3960 360 -3900 376
rect 2640 404 2700 420
rect 2640 376 2656 404
rect 2684 376 2700 404
rect 2640 360 2700 376
rect 2880 404 2940 420
rect 2880 376 2896 404
rect 2924 376 2940 404
rect 2880 360 2940 376
rect 4440 404 4500 420
rect 4440 376 4456 404
rect 4484 376 4500 404
rect 4440 360 4500 376
rect 4680 404 4740 420
rect 4680 376 4696 404
rect 4724 376 4740 404
rect 4680 360 4740 376
rect 5040 404 5100 420
rect 5040 376 5056 404
rect 5084 376 5100 404
rect 5040 360 5100 376
rect 5280 404 5340 420
rect 5280 376 5296 404
rect 5324 376 5340 404
rect 5280 360 5340 376
rect 6840 404 6900 420
rect 6840 376 6856 404
rect 6884 376 6900 404
rect 6840 360 6900 376
rect 7080 404 7140 420
rect 7080 376 7096 404
rect 7124 376 7140 404
rect 7080 360 7140 376
rect 13680 404 13740 420
rect 13680 376 13696 404
rect 13724 376 13740 404
rect 13680 360 13740 376
rect 14280 404 14340 420
rect 14280 376 14296 404
rect 14324 376 14340 404
rect 14280 360 14340 376
rect -5520 145 -5160 180
rect -5520 65 -5504 145
rect -5476 65 -5264 145
rect -5236 65 -5160 145
rect -5520 30 -5160 65
rect -2040 160 -1980 180
rect -2040 80 -2024 160
rect -1996 80 -1980 160
rect -2040 60 -1980 80
rect -960 160 -900 180
rect -960 80 -944 160
rect -916 80 -900 160
rect -960 60 -900 80
rect 2160 160 2220 180
rect 2160 80 2176 160
rect 2204 80 2220 160
rect 2160 60 2220 80
rect 2760 160 2820 180
rect 2760 80 2776 160
rect 2804 80 2820 160
rect 2760 60 2820 80
rect 4560 160 4620 180
rect 4560 80 4576 160
rect 4604 80 4620 160
rect 4560 60 4620 80
rect 5160 160 5220 180
rect 5160 80 5176 160
rect 5204 80 5220 160
rect 5160 60 5220 80
rect 6960 160 7020 180
rect 6960 80 6976 160
rect 7004 80 7020 160
rect 6960 60 7020 80
rect 7560 160 7620 180
rect 7560 80 7576 160
rect 7604 80 7620 160
rect 7560 60 7620 80
rect 10680 160 10740 180
rect 10680 80 10696 160
rect 10724 80 10740 160
rect 10680 60 10740 80
rect 11760 160 11820 180
rect 11760 80 11776 160
rect 11804 80 11820 160
rect 11760 60 11820 80
rect -5520 -16 -5160 0
rect -5520 -44 -5384 -16
rect -5356 -44 -5160 -16
rect -5520 -60 -5160 -44
rect -3720 -16 -3660 0
rect -3720 -44 -3704 -16
rect -3676 -44 -3660 -16
rect -3720 -60 -3660 -44
rect -3240 -16 -3180 0
rect -3240 -44 -3224 -16
rect -3196 -44 -3180 -16
rect -3240 -60 -3180 -44
rect -2760 -16 -2700 0
rect -2760 -44 -2744 -16
rect -2716 -44 -2700 -16
rect -2760 -60 -2700 -44
rect -2640 -16 -2580 0
rect -2640 -44 -2624 -16
rect -2596 -44 -2580 -16
rect -2640 -60 -2580 -44
rect -2160 -16 -2100 0
rect -2160 -44 -2144 -16
rect -2116 -44 -2100 -16
rect -2160 -60 -2100 -44
rect -1920 -16 -1860 0
rect -1920 -44 -1904 -16
rect -1876 -44 -1860 -16
rect -1920 -60 -1860 -44
rect 360 -16 420 0
rect 360 -44 376 -16
rect 404 -44 420 -16
rect 360 -60 420 -44
rect 2040 -16 2100 0
rect 2040 -44 2056 -16
rect 2084 -44 2100 -16
rect 2040 -60 2100 -44
rect 2280 -16 2340 0
rect 2280 -44 2296 -16
rect 2324 -44 2340 -16
rect 2280 -60 2340 -44
rect 7440 -16 7500 0
rect 7440 -44 7456 -16
rect 7484 -44 7500 -16
rect 7440 -60 7500 -44
rect 7680 -16 7740 0
rect 7680 -44 7696 -16
rect 7724 -44 7740 -16
rect 7680 -60 7740 -44
rect 9360 -16 9420 0
rect 9360 -44 9376 -16
rect 9404 -44 9420 -16
rect 9360 -60 9420 -44
rect 11640 -16 11700 0
rect 11640 -44 11656 -16
rect 11684 -44 11700 -16
rect 11640 -60 11700 -44
rect 11880 -16 11940 0
rect 11880 -44 11896 -16
rect 11924 -44 11940 -16
rect 11880 -60 11940 -44
rect 12360 -16 12420 0
rect 12360 -44 12376 -16
rect 12404 -44 12420 -16
rect 12360 -60 12420 -44
rect 12480 -16 12540 0
rect 12480 -44 12496 -16
rect 12524 -44 12540 -16
rect 12480 -60 12540 -44
rect 12960 -16 13020 0
rect 12960 -44 12976 -16
rect 13004 -44 13020 -16
rect 12960 -60 13020 -44
rect 13440 -16 13500 0
rect 13440 -44 13456 -16
rect 13484 -44 13500 -16
rect 13440 -60 13500 -44
rect -5520 -125 -5160 -90
rect -5520 -205 -5504 -125
rect -5476 -205 -5264 -125
rect -5236 -205 -5160 -125
rect -5520 -240 -5160 -205
rect -2040 -140 -1980 -120
rect -2040 -220 -2024 -140
rect -1996 -220 -1980 -140
rect -2040 -240 -1980 -220
rect -960 -140 -900 -120
rect -960 -220 -944 -140
rect -916 -220 -900 -140
rect -960 -240 -900 -220
rect 2160 -140 2220 -120
rect 2160 -220 2176 -140
rect 2204 -220 2220 -140
rect 2160 -240 2220 -220
rect 2760 -140 2820 -120
rect 2760 -220 2776 -140
rect 2804 -220 2820 -140
rect 2760 -240 2820 -220
rect 4560 -140 4620 -120
rect 4560 -220 4576 -140
rect 4604 -220 4620 -140
rect 4560 -240 4620 -220
rect 5160 -140 5220 -120
rect 5160 -220 5176 -140
rect 5204 -220 5220 -140
rect 5160 -240 5220 -220
rect 6960 -140 7020 -120
rect 6960 -220 6976 -140
rect 7004 -220 7020 -140
rect 6960 -240 7020 -220
rect 7560 -140 7620 -120
rect 7560 -220 7576 -140
rect 7604 -220 7620 -140
rect 7560 -240 7620 -220
rect 10680 -140 10740 -120
rect 10680 -220 10696 -140
rect 10724 -220 10740 -140
rect 10680 -240 10740 -220
rect 11760 -140 11820 -120
rect 11760 -220 11776 -140
rect 11804 -220 11820 -140
rect 11760 -240 11820 -220
rect -5220 -840 -5160 -540
<< via3 >>
rect -5504 1385 -5476 1465
rect -5264 1385 -5236 1465
rect -104 1400 -76 1480
rect 9856 1400 9884 1480
rect -5384 1276 -5356 1304
rect -4304 1276 -4276 1304
rect -3344 1276 -3316 1304
rect -1544 1276 -1516 1304
rect -1304 1276 -1276 1304
rect 1456 1276 1484 1304
rect 1696 1276 1724 1304
rect 8056 1276 8084 1304
rect 8296 1276 8324 1304
rect 11056 1276 11084 1304
rect 11296 1276 11324 1304
rect 13096 1276 13124 1304
rect 14056 1276 14084 1304
rect -5504 1115 -5476 1195
rect -5264 1115 -5236 1195
rect -104 1100 -76 1180
rect 9856 1100 9884 1180
rect -3104 856 -3076 884
rect -2504 856 -2476 884
rect 3256 856 3284 884
rect 3496 856 3524 884
rect 3856 856 3884 884
rect 4096 856 4124 884
rect 5656 856 5684 884
rect 5896 856 5924 884
rect 6256 856 6284 884
rect 6496 856 6524 884
rect 12256 856 12284 884
rect 12856 856 12884 884
rect -704 616 -676 644
rect -344 616 -316 644
rect 256 616 284 644
rect 496 616 524 644
rect 856 616 884 644
rect 1096 616 1124 644
rect 8656 616 8684 644
rect 8896 616 8924 644
rect 9256 616 9284 644
rect 9496 616 9524 644
rect 10096 616 10124 644
rect 10456 616 10484 644
rect -4544 376 -4516 404
rect -3944 376 -3916 404
rect 2656 376 2684 404
rect 2896 376 2924 404
rect 4456 376 4484 404
rect 4696 376 4724 404
rect 5056 376 5084 404
rect 5296 376 5324 404
rect 6856 376 6884 404
rect 7096 376 7124 404
rect 13696 376 13724 404
rect 14296 376 14324 404
rect -5504 65 -5476 145
rect -5264 65 -5236 145
rect -944 80 -916 160
rect 10696 80 10724 160
rect -5384 -44 -5356 -16
rect -3704 -44 -3676 -16
rect -2744 -44 -2716 -16
rect -2144 -44 -2116 -16
rect -1904 -44 -1876 -16
rect 2056 -44 2084 -16
rect 2296 -44 2324 -16
rect 7456 -44 7484 -16
rect 7696 -44 7724 -16
rect 11656 -44 11684 -16
rect 11896 -44 11924 -16
rect 12496 -44 12524 -16
rect 13456 -44 13484 -16
rect -5504 -205 -5476 -125
rect -5264 -205 -5236 -125
rect -944 -220 -916 -140
rect 10696 -220 10724 -140
<< metal4 >>
rect -5160 4200 14940 4260
rect -5520 3464 -5460 3540
rect -5520 3436 -5504 3464
rect -5476 3436 -5460 3464
rect -5520 3224 -5460 3436
rect -5520 3196 -5504 3224
rect -5476 3196 -5460 3224
rect -5520 1465 -5460 3196
rect -5520 1385 -5504 1465
rect -5476 1385 -5460 1465
rect -5520 1195 -5460 1385
rect -5520 1115 -5504 1195
rect -5476 1115 -5460 1195
rect -5520 1080 -5460 1115
rect -5400 3344 -5340 3540
rect -5400 3316 -5384 3344
rect -5356 3316 -5340 3344
rect -5400 1304 -5340 3316
rect -5400 1276 -5384 1304
rect -5356 1276 -5340 1304
rect -5400 1080 -5340 1276
rect -5280 3464 -5220 3540
rect -5280 3436 -5264 3464
rect -5236 3436 -5220 3464
rect -5280 3224 -5220 3436
rect -5160 3480 -5100 4200
rect 14880 3480 14940 4200
rect -5160 3344 14940 3480
rect -5160 3316 -5082 3344
rect 14862 3316 14940 3344
rect -5160 3300 14940 3316
rect -5280 3196 -5264 3224
rect -5236 3196 -5220 3224
rect -5280 1465 -5220 3196
rect -5280 1385 -5264 1465
rect -5236 1385 -5220 1465
rect -5280 1195 -5220 1385
rect -120 1480 -60 1500
rect -120 1400 -104 1480
rect -76 1400 -60 1480
rect -120 1380 -60 1400
rect 9840 1480 9900 1500
rect 9840 1400 9856 1480
rect 9884 1400 9900 1480
rect 9840 1380 9900 1400
rect -4320 1304 -4260 1320
rect -4320 1276 -4304 1304
rect -4276 1276 -4260 1304
rect -4320 1260 -4260 1276
rect -3360 1304 -3300 1320
rect -3360 1276 -3344 1304
rect -3316 1276 -3300 1304
rect -3360 1260 -3300 1276
rect -1560 1304 -1500 1320
rect -1560 1276 -1544 1304
rect -1516 1276 -1500 1304
rect -1560 1260 -1500 1276
rect -1320 1304 -1260 1320
rect -1320 1276 -1304 1304
rect -1276 1276 -1260 1304
rect -1320 1260 -1260 1276
rect 1440 1304 1500 1320
rect 1440 1276 1456 1304
rect 1484 1276 1500 1304
rect 1440 1260 1500 1276
rect 1680 1304 1740 1320
rect 1680 1276 1696 1304
rect 1724 1276 1740 1304
rect 1680 1260 1740 1276
rect 8040 1304 8100 1320
rect 8040 1276 8056 1304
rect 8084 1276 8100 1304
rect 8040 1260 8100 1276
rect 8280 1304 8340 1320
rect 8280 1276 8296 1304
rect 8324 1276 8340 1304
rect 8280 1260 8340 1276
rect 11040 1304 11100 1320
rect 11040 1276 11056 1304
rect 11084 1276 11100 1304
rect 11040 1260 11100 1276
rect 11280 1304 11340 1320
rect 11280 1276 11296 1304
rect 11324 1276 11340 1304
rect 11280 1260 11340 1276
rect 13080 1304 13140 1320
rect 13080 1276 13096 1304
rect 13124 1276 13140 1304
rect 13080 1260 13140 1276
rect 14040 1304 14100 1320
rect 14040 1276 14056 1304
rect 14084 1276 14100 1304
rect 14040 1260 14100 1276
rect -5280 1115 -5264 1195
rect -5236 1115 -5220 1195
rect -5280 1080 -5220 1115
rect -120 1180 -60 1200
rect -120 1100 -104 1180
rect -76 1100 -60 1180
rect -120 1080 -60 1100
rect 9840 1180 9900 1200
rect 9840 1100 9856 1180
rect 9884 1100 9900 1180
rect 9840 1080 9900 1100
rect -3120 884 -3060 900
rect -3120 856 -3104 884
rect -3076 856 -3060 884
rect -3120 840 -3060 856
rect -2520 884 -2460 900
rect -2520 856 -2504 884
rect -2476 856 -2460 884
rect -2520 840 -2460 856
rect 3240 884 3300 900
rect 3240 856 3256 884
rect 3284 856 3300 884
rect 3240 840 3300 856
rect 3480 884 3540 900
rect 3480 856 3496 884
rect 3524 856 3540 884
rect 3480 840 3540 856
rect 3840 884 3900 900
rect 3840 856 3856 884
rect 3884 856 3900 884
rect 3840 840 3900 856
rect 4080 884 4140 900
rect 4080 856 4096 884
rect 4124 856 4140 884
rect 4080 840 4140 856
rect 5640 884 5700 900
rect 5640 856 5656 884
rect 5684 856 5700 884
rect 5640 840 5700 856
rect 5880 884 5940 900
rect 5880 856 5896 884
rect 5924 856 5940 884
rect 5880 840 5940 856
rect 6240 884 6300 900
rect 6240 856 6256 884
rect 6284 856 6300 884
rect 6240 840 6300 856
rect 6480 884 6540 900
rect 6480 856 6496 884
rect 6524 856 6540 884
rect 6480 840 6540 856
rect 12240 884 12300 900
rect 12240 856 12256 884
rect 12284 856 12300 884
rect 12240 840 12300 856
rect 12840 884 12900 900
rect 12840 856 12856 884
rect 12884 856 12900 884
rect 12840 840 12900 856
rect -720 644 -660 660
rect -720 616 -704 644
rect -676 616 -660 644
rect -720 600 -660 616
rect -360 644 -300 660
rect -360 616 -344 644
rect -316 616 -300 644
rect -360 600 -300 616
rect 240 644 300 660
rect 240 616 256 644
rect 284 616 300 644
rect 240 600 300 616
rect 480 644 540 660
rect 480 616 496 644
rect 524 616 540 644
rect 480 600 540 616
rect 840 644 900 660
rect 840 616 856 644
rect 884 616 900 644
rect 840 600 900 616
rect 1080 644 1140 660
rect 1080 616 1096 644
rect 1124 616 1140 644
rect 1080 600 1140 616
rect 8640 644 8700 660
rect 8640 616 8656 644
rect 8684 616 8700 644
rect 8640 600 8700 616
rect 8880 644 8940 660
rect 8880 616 8896 644
rect 8924 616 8940 644
rect 8880 600 8940 616
rect 9240 644 9300 660
rect 9240 616 9256 644
rect 9284 616 9300 644
rect 9240 600 9300 616
rect 9480 644 9540 660
rect 9480 616 9496 644
rect 9524 616 9540 644
rect 9480 600 9540 616
rect 10080 644 10140 660
rect 10080 616 10096 644
rect 10124 616 10140 644
rect 10080 600 10140 616
rect 10440 644 10500 660
rect 10440 616 10456 644
rect 10484 616 10500 644
rect 10440 600 10500 616
rect -4560 404 -4500 420
rect -4560 376 -4544 404
rect -4516 376 -4500 404
rect -4560 360 -4500 376
rect -3960 404 -3900 420
rect -3960 376 -3944 404
rect -3916 376 -3900 404
rect -3960 360 -3900 376
rect 2640 404 2700 420
rect 2640 376 2656 404
rect 2684 376 2700 404
rect 2640 360 2700 376
rect 2880 404 2940 420
rect 2880 376 2896 404
rect 2924 376 2940 404
rect 2880 360 2940 376
rect 4440 404 4500 420
rect 4440 376 4456 404
rect 4484 376 4500 404
rect 4440 360 4500 376
rect 4680 404 4740 420
rect 4680 376 4696 404
rect 4724 376 4740 404
rect 4680 360 4740 376
rect 5040 404 5100 420
rect 5040 376 5056 404
rect 5084 376 5100 404
rect 5040 360 5100 376
rect 5280 404 5340 420
rect 5280 376 5296 404
rect 5324 376 5340 404
rect 5280 360 5340 376
rect 6840 404 6900 420
rect 6840 376 6856 404
rect 6884 376 6900 404
rect 6840 360 6900 376
rect 7080 404 7140 420
rect 7080 376 7096 404
rect 7124 376 7140 404
rect 7080 360 7140 376
rect 13680 404 13740 420
rect 13680 376 13696 404
rect 13724 376 13740 404
rect 13680 360 13740 376
rect 14280 404 14340 420
rect 14280 376 14296 404
rect 14324 376 14340 404
rect 14280 360 14340 376
rect -5520 145 -5460 180
rect -5520 65 -5504 145
rect -5476 65 -5460 145
rect -5520 -125 -5460 65
rect -5520 -205 -5504 -125
rect -5476 -205 -5460 -125
rect -5520 -916 -5460 -205
rect -5520 -944 -5504 -916
rect -5476 -944 -5460 -916
rect -5520 -1156 -5460 -944
rect -5520 -1184 -5504 -1156
rect -5476 -1184 -5460 -1156
rect -5520 -1260 -5460 -1184
rect -5400 -16 -5340 180
rect -5400 -44 -5384 -16
rect -5356 -44 -5340 -16
rect -5400 -1036 -5340 -44
rect -5400 -1064 -5384 -1036
rect -5356 -1064 -5340 -1036
rect -5400 -1260 -5340 -1064
rect -5280 145 -5220 180
rect -5280 65 -5264 145
rect -5236 65 -5220 145
rect -5280 -125 -5220 65
rect -960 160 -900 180
rect -960 80 -944 160
rect -916 80 -900 160
rect -960 60 -900 80
rect 10680 160 10740 180
rect 10680 80 10696 160
rect 10724 80 10740 160
rect 10680 60 10740 80
rect -3720 -16 -3660 0
rect -3720 -44 -3704 -16
rect -3676 -44 -3660 -16
rect -3720 -60 -3660 -44
rect -2760 -16 -2700 0
rect -2760 -44 -2744 -16
rect -2716 -44 -2700 -16
rect -2760 -60 -2700 -44
rect -2160 -16 -2100 0
rect -2160 -44 -2144 -16
rect -2116 -44 -2100 -16
rect -2160 -60 -2100 -44
rect -1920 -16 -1860 0
rect -1920 -44 -1904 -16
rect -1876 -44 -1860 -16
rect -1920 -60 -1860 -44
rect 2040 -16 2100 0
rect 2040 -44 2056 -16
rect 2084 -44 2100 -16
rect 2040 -60 2100 -44
rect 2280 -16 2340 0
rect 2280 -44 2296 -16
rect 2324 -44 2340 -16
rect 2280 -60 2340 -44
rect 7440 -16 7500 0
rect 7440 -44 7456 -16
rect 7484 -44 7500 -16
rect 7440 -60 7500 -44
rect 7680 -16 7740 0
rect 7680 -44 7696 -16
rect 7724 -44 7740 -16
rect 7680 -60 7740 -44
rect 11640 -16 11700 0
rect 11640 -44 11656 -16
rect 11684 -44 11700 -16
rect 11640 -60 11700 -44
rect 11880 -16 11940 0
rect 11880 -44 11896 -16
rect 11924 -44 11940 -16
rect 11880 -60 11940 -44
rect 12480 -16 12540 0
rect 12480 -44 12496 -16
rect 12524 -44 12540 -16
rect 12480 -60 12540 -44
rect 13440 -16 13500 0
rect 13440 -44 13456 -16
rect 13484 -44 13500 -16
rect 13440 -60 13500 -44
rect -5280 -205 -5264 -125
rect -5236 -205 -5220 -125
rect -5280 -916 -5220 -205
rect -960 -140 -900 -120
rect -960 -220 -944 -140
rect -916 -220 -900 -140
rect -960 -240 -900 -220
rect 10680 -140 10740 -120
rect 10680 -220 10696 -140
rect 10724 -220 10740 -140
rect 10680 -240 10740 -220
rect -5280 -944 -5264 -916
rect -5236 -944 -5220 -916
rect -5280 -1156 -5220 -944
rect -5280 -1184 -5264 -1156
rect -5236 -1184 -5220 -1156
rect -5280 -1260 -5220 -1184
rect -5160 -1036 14940 -1020
rect -5160 -1064 -5082 -1036
rect 14862 -1064 14940 -1036
rect -5160 -1200 14940 -1064
rect -5160 -1920 -5100 -1200
rect 14880 -1920 14940 -1200
rect -5160 -1980 14940 -1920
<< via4 >>
rect -5504 3436 -5476 3464
rect -5504 3196 -5476 3224
rect -5384 3316 -5356 3344
rect -5264 3436 -5236 3464
rect -5082 3316 14862 3344
rect -5264 3196 -5236 3224
rect -5504 -944 -5476 -916
rect -5504 -1184 -5476 -1156
rect -5384 -1064 -5356 -1036
rect -5264 -944 -5236 -916
rect -5264 -1184 -5236 -1156
rect -5082 -1064 14862 -1036
<< metal5 >>
rect -5160 3962 14940 4260
rect -5160 3538 -5042 3962
rect -4618 3538 14940 3962
rect -5160 3480 14940 3538
rect -5580 3464 14940 3480
rect -5580 3436 -5504 3464
rect -5476 3436 -5264 3464
rect -5236 3436 14940 3464
rect -5580 3420 14940 3436
rect -5580 3344 14940 3360
rect -5580 3316 -5384 3344
rect -5356 3316 -5082 3344
rect 14862 3316 14940 3344
rect -5580 3300 14940 3316
rect -5580 3224 14940 3240
rect -5580 3196 -5504 3224
rect -5476 3196 -5264 3224
rect -5236 3196 14940 3224
rect -5580 3180 14940 3196
rect -5580 -916 14940 -900
rect -5580 -944 -5504 -916
rect -5476 -944 -5264 -916
rect -5236 -944 14940 -916
rect -5580 -960 14940 -944
rect -5580 -1036 14940 -1020
rect -5580 -1064 -5384 -1036
rect -5356 -1064 -5082 -1036
rect 14862 -1064 14940 -1036
rect -5580 -1080 14940 -1064
rect -5580 -1156 14940 -1140
rect -5580 -1184 -5504 -1156
rect -5476 -1184 -5264 -1156
rect -5236 -1184 14940 -1156
rect -5580 -1200 14940 -1184
rect -5160 -1258 14940 -1200
rect -5160 -1682 -5042 -1258
rect -4618 -1682 14940 -1258
rect -5160 -1980 14940 -1682
use nautavieru_cell#0  nautavieru_cell_0
timestamp 1665184495
transform -1 0 10920 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_1
timestamp 1665184495
transform -1 0 10320 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_2
timestamp 1665184495
transform -1 0 9120 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_3
timestamp 1665184495
transform -1 0 9720 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_4
timestamp 1665184495
transform -1 0 8520 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_5
timestamp 1665184495
transform -1 0 7920 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_6
timestamp 1665184495
transform -1 0 7320 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_7
timestamp 1665184495
transform -1 0 6720 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_8
timestamp 1665184495
transform -1 0 6120 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_9
timestamp 1665184495
transform -1 0 5520 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_10
timestamp 1665184495
transform -1 0 4920 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_11
timestamp 1665184495
transform -1 0 4320 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_12
timestamp 1665184495
transform -1 0 3720 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_13
timestamp 1665184495
transform -1 0 3120 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_14
timestamp 1665184495
transform -1 0 2520 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_15
timestamp 1665184495
transform -1 0 1920 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_16
timestamp 1665184495
transform 1 0 7860 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_17
timestamp 1665184495
transform 1 0 7260 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_18
timestamp 1665184495
transform 1 0 6660 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_19
timestamp 1665184495
transform 1 0 6060 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_20
timestamp 1665184495
transform 1 0 5460 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_21
timestamp 1665184495
transform 1 0 4860 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_22
timestamp 1665184495
transform 1 0 4260 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_23
timestamp 1665184495
transform 1 0 3660 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_24
timestamp 1665184495
transform 1 0 3060 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_25
timestamp 1665184495
transform 1 0 2460 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_26
timestamp 1665184495
transform 1 0 1860 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_27
timestamp 1665184495
transform 1 0 1260 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_28
timestamp 1665184495
transform 1 0 660 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_29
timestamp 1665184495
transform 1 0 60 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_30
timestamp 1665184495
transform 1 0 -540 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_cell#0  nautavieru_cell_31
timestamp 1665184495
transform 1 0 -1140 0 1 -180
box -3600 -660 -2940 3300
use nautavieru_edge#0  nautavieru_edge_0
timestamp 1665184495
transform -1 0 11160 0 1 -180
box -3780 -660 -3300 3300
use nautavieru_edge#0  nautavieru_edge_1
timestamp 1665184495
transform 1 0 -1380 0 1 -180
box -3780 -660 -3300 3300
<< labels >>
rlabel metal3 s -5190 -30 -5190 -30 4 xp
rlabel metal3 s -5190 1290 -5190 1290 4 xm
rlabel metal3 s -5190 630 -5190 630 4 x
rlabel metal3 s -5220 360 -5160 420 4 ip
port 1 nsew
rlabel metal3 s -5220 840 -5160 900 4 im
port 2 nsew
rlabel metal3 s -5220 1440 -5160 1500 4 op
port 3 nsew
rlabel metal3 s -5220 -240 -5160 -180 4 om
port 4 nsew
rlabel metal3 s -5220 2700 -5160 3000 4 vdd
port 5 nsew
rlabel metal3 s -5220 2340 -5160 2400 4 gp
port 6 nsew
rlabel metal3 s -5220 1680 -5160 1740 4 bp
port 7 nsew
rlabel metal3 s -5220 2460 -5160 2520 4 vreg
port 8 nsew
rlabel metal3 s -5220 -840 -5160 -540 4 gnd
port 9 nsew
<< end >>
