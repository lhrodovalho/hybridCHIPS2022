magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7200 5220 -5880 6420
rect -7200 3660 -5880 4980
<< nmos >>
rect -6960 -1080 -6840 -720
rect -6720 -1080 -6600 -720
rect -6480 -1080 -6360 -720
rect -6240 -1080 -6120 -720
<< pmos >>
rect -6960 4200 -6840 4500
rect -6720 4200 -6600 4500
rect -6480 4200 -6360 4500
rect -6240 4200 -6120 4500
<< mvpmos >>
rect -6960 5760 -6840 6120
rect -6720 5760 -6600 6120
rect -6480 5760 -6360 6120
rect -6240 5760 -6120 6120
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -757 -6480 -720
rect -6600 -803 -6563 -757
rect -6517 -803 -6480 -757
rect -6600 -877 -6480 -803
rect -6600 -923 -6563 -877
rect -6517 -923 -6480 -877
rect -6600 -997 -6480 -923
rect -6600 -1043 -6563 -997
rect -6517 -1043 -6480 -997
rect -6600 -1080 -6480 -1043
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -757 -6000 -720
rect -6120 -803 -6083 -757
rect -6037 -803 -6000 -757
rect -6120 -877 -6000 -803
rect -6120 -923 -6083 -877
rect -6037 -923 -6000 -877
rect -6120 -997 -6000 -923
rect -6120 -1043 -6083 -997
rect -6037 -1043 -6000 -997
rect -6120 -1080 -6000 -1043
<< pdiff >>
rect -7080 4403 -6960 4500
rect -7080 4357 -7043 4403
rect -6997 4357 -6960 4403
rect -7080 4283 -6960 4357
rect -7080 4237 -7043 4283
rect -6997 4237 -6960 4283
rect -7080 4200 -6960 4237
rect -6840 4403 -6720 4500
rect -6840 4357 -6803 4403
rect -6757 4357 -6720 4403
rect -6840 4283 -6720 4357
rect -6840 4237 -6803 4283
rect -6757 4237 -6720 4283
rect -6840 4200 -6720 4237
rect -6600 4403 -6480 4500
rect -6600 4357 -6563 4403
rect -6517 4357 -6480 4403
rect -6600 4283 -6480 4357
rect -6600 4237 -6563 4283
rect -6517 4237 -6480 4283
rect -6600 4200 -6480 4237
rect -6360 4403 -6240 4500
rect -6360 4357 -6323 4403
rect -6277 4357 -6240 4403
rect -6360 4283 -6240 4357
rect -6360 4237 -6323 4283
rect -6277 4237 -6240 4283
rect -6360 4200 -6240 4237
rect -6120 4403 -6000 4500
rect -6120 4357 -6083 4403
rect -6037 4357 -6000 4403
rect -6120 4283 -6000 4357
rect -6120 4237 -6083 4283
rect -6037 4237 -6000 4283
rect -6120 4200 -6000 4237
<< mvpdiff >>
rect -7080 6083 -6960 6120
rect -7080 6037 -7043 6083
rect -6997 6037 -6960 6083
rect -7080 5963 -6960 6037
rect -7080 5917 -7043 5963
rect -6997 5917 -6960 5963
rect -7080 5843 -6960 5917
rect -7080 5797 -7043 5843
rect -6997 5797 -6960 5843
rect -7080 5760 -6960 5797
rect -6840 6083 -6720 6120
rect -6840 6037 -6803 6083
rect -6757 6037 -6720 6083
rect -6840 5963 -6720 6037
rect -6840 5917 -6803 5963
rect -6757 5917 -6720 5963
rect -6840 5843 -6720 5917
rect -6840 5797 -6803 5843
rect -6757 5797 -6720 5843
rect -6840 5760 -6720 5797
rect -6600 6083 -6480 6120
rect -6600 6037 -6563 6083
rect -6517 6037 -6480 6083
rect -6600 5963 -6480 6037
rect -6600 5917 -6563 5963
rect -6517 5917 -6480 5963
rect -6600 5843 -6480 5917
rect -6600 5797 -6563 5843
rect -6517 5797 -6480 5843
rect -6600 5760 -6480 5797
rect -6360 6083 -6240 6120
rect -6360 6037 -6323 6083
rect -6277 6037 -6240 6083
rect -6360 5963 -6240 6037
rect -6360 5917 -6323 5963
rect -6277 5917 -6240 5963
rect -6360 5843 -6240 5917
rect -6360 5797 -6323 5843
rect -6277 5797 -6240 5843
rect -6360 5760 -6240 5797
rect -6120 6083 -6000 6120
rect -6120 6037 -6083 6083
rect -6037 6037 -6000 6083
rect -6120 5963 -6000 6037
rect -6120 5917 -6083 5963
rect -6037 5917 -6000 5963
rect -6120 5843 -6000 5917
rect -6120 5797 -6083 5843
rect -6037 5797 -6000 5843
rect -6120 5760 -6000 5797
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
rect -6563 -803 -6517 -757
rect -6563 -923 -6517 -877
rect -6563 -1043 -6517 -997
rect -6323 -803 -6277 -757
rect -6323 -923 -6277 -877
rect -6323 -1043 -6277 -997
rect -6083 -803 -6037 -757
rect -6083 -923 -6037 -877
rect -6083 -1043 -6037 -997
<< pdiffc >>
rect -7043 4357 -6997 4403
rect -7043 4237 -6997 4283
rect -6803 4357 -6757 4403
rect -6803 4237 -6757 4283
rect -6563 4357 -6517 4403
rect -6563 4237 -6517 4283
rect -6323 4357 -6277 4403
rect -6323 4237 -6277 4283
rect -6083 4357 -6037 4403
rect -6083 4237 -6037 4283
<< mvpdiffc >>
rect -7043 6037 -6997 6083
rect -7043 5917 -6997 5963
rect -7043 5797 -6997 5843
rect -6803 6037 -6757 6083
rect -6803 5917 -6757 5963
rect -6803 5797 -6757 5843
rect -6563 6037 -6517 6083
rect -6563 5917 -6517 5963
rect -6563 5797 -6517 5843
rect -6323 6037 -6277 6083
rect -6323 5917 -6277 5963
rect -6323 5797 -6277 5843
rect -6083 6037 -6037 6083
rect -6083 5917 -6037 5963
rect -6083 5797 -6037 5843
<< psubdiff >>
rect -7200 6563 -5880 6600
rect -7200 6517 -7163 6563
rect -7117 6517 -7043 6563
rect -6997 6517 -6923 6563
rect -6877 6517 -6803 6563
rect -6757 6517 -6683 6563
rect -6637 6517 -6563 6563
rect -6517 6517 -6443 6563
rect -6397 6517 -6323 6563
rect -6277 6517 -6203 6563
rect -6157 6517 -6083 6563
rect -6037 6517 -5963 6563
rect -5917 6517 -5880 6563
rect -7200 6480 -5880 6517
rect -7200 5123 -5880 5160
rect -7200 5077 -7163 5123
rect -7117 5077 -7043 5123
rect -6997 5077 -6923 5123
rect -6877 5077 -6803 5123
rect -6757 5077 -6683 5123
rect -6637 5077 -6563 5123
rect -6517 5077 -6443 5123
rect -6397 5077 -6323 5123
rect -6277 5077 -6203 5123
rect -6157 5077 -6083 5123
rect -6037 5077 -5963 5123
rect -5917 5077 -5880 5123
rect -7200 5040 -5880 5077
rect -7200 3563 -5880 3600
rect -7200 3517 -7163 3563
rect -7117 3517 -7043 3563
rect -6997 3517 -6923 3563
rect -6877 3517 -6803 3563
rect -6757 3517 -6683 3563
rect -6637 3517 -6563 3563
rect -6517 3517 -6443 3563
rect -6397 3517 -6323 3563
rect -6277 3517 -6203 3563
rect -6157 3517 -6083 3563
rect -6037 3517 -5963 3563
rect -5917 3517 -5880 3563
rect -7200 3480 -5880 3517
rect -7200 2603 -5880 2640
rect -7200 2557 -7163 2603
rect -7117 2557 -7043 2603
rect -6997 2557 -6923 2603
rect -6877 2557 -6803 2603
rect -6757 2557 -6683 2603
rect -6637 2557 -6563 2603
rect -6517 2557 -6443 2603
rect -6397 2557 -6323 2603
rect -6277 2557 -6203 2603
rect -6157 2557 -6083 2603
rect -6037 2557 -5963 2603
rect -5917 2557 -5880 2603
rect -7200 2520 -5880 2557
rect -7200 2123 -5880 2160
rect -7200 2077 -7163 2123
rect -7117 2077 -7043 2123
rect -6997 2077 -6923 2123
rect -6877 2077 -6803 2123
rect -6757 2077 -6683 2123
rect -6637 2077 -6563 2123
rect -6517 2077 -6443 2123
rect -6397 2077 -6323 2123
rect -6277 2077 -6203 2123
rect -6157 2077 -6083 2123
rect -6037 2077 -5963 2123
rect -5917 2077 -5880 2123
rect -7200 2040 -5880 2077
rect -7200 1643 -5880 1680
rect -7200 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6563 1643
rect -6517 1597 -6443 1643
rect -6397 1597 -6323 1643
rect -6277 1597 -6203 1643
rect -6157 1597 -6083 1643
rect -6037 1597 -5963 1643
rect -5917 1597 -5880 1643
rect -7200 1560 -5880 1597
rect -7200 1163 -5880 1200
rect -7200 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6563 1163
rect -6517 1117 -6443 1163
rect -6397 1117 -6323 1163
rect -6277 1117 -6203 1163
rect -6157 1117 -6083 1163
rect -6037 1117 -5963 1163
rect -5917 1117 -5880 1163
rect -7200 1080 -5880 1117
rect -7200 683 -5880 720
rect -7200 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6563 683
rect -6517 637 -6443 683
rect -6397 637 -6323 683
rect -6277 637 -6203 683
rect -6157 637 -6083 683
rect -6037 637 -5963 683
rect -5917 637 -5880 683
rect -7200 600 -5880 637
rect -7200 -277 -5880 -240
rect -7200 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6083 -277
rect -6037 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -360 -5880 -323
rect -7200 -1237 -5880 -1200
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6083 -1237
rect -6037 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1320 -5880 -1283
<< nsubdiff >>
rect -7080 4883 -6000 4920
rect -7080 4837 -7043 4883
rect -6997 4837 -6923 4883
rect -6877 4837 -6803 4883
rect -6757 4837 -6683 4883
rect -6637 4837 -6563 4883
rect -6517 4837 -6443 4883
rect -6397 4837 -6323 4883
rect -6277 4837 -6203 4883
rect -6157 4837 -6083 4883
rect -6037 4837 -6000 4883
rect -7080 4800 -6000 4837
rect -7080 3803 -6000 3840
rect -7080 3757 -7043 3803
rect -6997 3757 -6923 3803
rect -6877 3757 -6803 3803
rect -6757 3757 -6683 3803
rect -6637 3757 -6563 3803
rect -6517 3757 -6443 3803
rect -6397 3757 -6323 3803
rect -6277 3757 -6203 3803
rect -6157 3757 -6083 3803
rect -6037 3757 -6000 3803
rect -7080 3720 -6000 3757
<< mvnsubdiff >>
rect -7080 6323 -6000 6360
rect -7080 6277 -7043 6323
rect -6997 6277 -6923 6323
rect -6877 6277 -6803 6323
rect -6757 6277 -6683 6323
rect -6637 6277 -6563 6323
rect -6517 6277 -6443 6323
rect -6397 6277 -6323 6323
rect -6277 6277 -6203 6323
rect -6157 6277 -6083 6323
rect -6037 6277 -6000 6323
rect -7080 6240 -6000 6277
rect -7080 5363 -6000 5400
rect -7080 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6683 5363
rect -6637 5317 -6563 5363
rect -6517 5317 -6443 5363
rect -6397 5317 -6323 5363
rect -6277 5317 -6203 5363
rect -6157 5317 -6083 5363
rect -6037 5317 -6000 5363
rect -7080 5280 -6000 5317
<< psubdiffcont >>
rect -7163 6517 -7117 6563
rect -7043 6517 -6997 6563
rect -6923 6517 -6877 6563
rect -6803 6517 -6757 6563
rect -6683 6517 -6637 6563
rect -6563 6517 -6517 6563
rect -6443 6517 -6397 6563
rect -6323 6517 -6277 6563
rect -6203 6517 -6157 6563
rect -6083 6517 -6037 6563
rect -5963 6517 -5917 6563
rect -7163 5077 -7117 5123
rect -7043 5077 -6997 5123
rect -6923 5077 -6877 5123
rect -6803 5077 -6757 5123
rect -6683 5077 -6637 5123
rect -6563 5077 -6517 5123
rect -6443 5077 -6397 5123
rect -6323 5077 -6277 5123
rect -6203 5077 -6157 5123
rect -6083 5077 -6037 5123
rect -5963 5077 -5917 5123
rect -7163 3517 -7117 3563
rect -7043 3517 -6997 3563
rect -6923 3517 -6877 3563
rect -6803 3517 -6757 3563
rect -6683 3517 -6637 3563
rect -6563 3517 -6517 3563
rect -6443 3517 -6397 3563
rect -6323 3517 -6277 3563
rect -6203 3517 -6157 3563
rect -6083 3517 -6037 3563
rect -5963 3517 -5917 3563
rect -7163 2557 -7117 2603
rect -7043 2557 -6997 2603
rect -6923 2557 -6877 2603
rect -6803 2557 -6757 2603
rect -6683 2557 -6637 2603
rect -6563 2557 -6517 2603
rect -6443 2557 -6397 2603
rect -6323 2557 -6277 2603
rect -6203 2557 -6157 2603
rect -6083 2557 -6037 2603
rect -5963 2557 -5917 2603
rect -7163 2077 -7117 2123
rect -7043 2077 -6997 2123
rect -6923 2077 -6877 2123
rect -6803 2077 -6757 2123
rect -6683 2077 -6637 2123
rect -6563 2077 -6517 2123
rect -6443 2077 -6397 2123
rect -6323 2077 -6277 2123
rect -6203 2077 -6157 2123
rect -6083 2077 -6037 2123
rect -5963 2077 -5917 2123
rect -7163 1597 -7117 1643
rect -7043 1597 -6997 1643
rect -6923 1597 -6877 1643
rect -6803 1597 -6757 1643
rect -6683 1597 -6637 1643
rect -6563 1597 -6517 1643
rect -6443 1597 -6397 1643
rect -6323 1597 -6277 1643
rect -6203 1597 -6157 1643
rect -6083 1597 -6037 1643
rect -5963 1597 -5917 1643
rect -7163 1117 -7117 1163
rect -7043 1117 -6997 1163
rect -6923 1117 -6877 1163
rect -6803 1117 -6757 1163
rect -6683 1117 -6637 1163
rect -6563 1117 -6517 1163
rect -6443 1117 -6397 1163
rect -6323 1117 -6277 1163
rect -6203 1117 -6157 1163
rect -6083 1117 -6037 1163
rect -5963 1117 -5917 1163
rect -7163 637 -7117 683
rect -7043 637 -6997 683
rect -6923 637 -6877 683
rect -6803 637 -6757 683
rect -6683 637 -6637 683
rect -6563 637 -6517 683
rect -6443 637 -6397 683
rect -6323 637 -6277 683
rect -6203 637 -6157 683
rect -6083 637 -6037 683
rect -5963 637 -5917 683
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -6563 -323 -6517 -277
rect -6443 -323 -6397 -277
rect -6323 -323 -6277 -277
rect -6203 -323 -6157 -277
rect -6083 -323 -6037 -277
rect -5963 -323 -5917 -277
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
rect -6563 -1283 -6517 -1237
rect -6443 -1283 -6397 -1237
rect -6323 -1283 -6277 -1237
rect -6203 -1283 -6157 -1237
rect -6083 -1283 -6037 -1237
rect -5963 -1283 -5917 -1237
<< nsubdiffcont >>
rect -7043 4837 -6997 4883
rect -6923 4837 -6877 4883
rect -6803 4837 -6757 4883
rect -6683 4837 -6637 4883
rect -6563 4837 -6517 4883
rect -6443 4837 -6397 4883
rect -6323 4837 -6277 4883
rect -6203 4837 -6157 4883
rect -6083 4837 -6037 4883
rect -7043 3757 -6997 3803
rect -6923 3757 -6877 3803
rect -6803 3757 -6757 3803
rect -6683 3757 -6637 3803
rect -6563 3757 -6517 3803
rect -6443 3757 -6397 3803
rect -6323 3757 -6277 3803
rect -6203 3757 -6157 3803
rect -6083 3757 -6037 3803
<< mvnsubdiffcont >>
rect -7043 6277 -6997 6323
rect -6923 6277 -6877 6323
rect -6803 6277 -6757 6323
rect -6683 6277 -6637 6323
rect -6563 6277 -6517 6323
rect -6443 6277 -6397 6323
rect -6323 6277 -6277 6323
rect -6203 6277 -6157 6323
rect -6083 6277 -6037 6323
rect -7043 5317 -6997 5363
rect -6923 5317 -6877 5363
rect -6803 5317 -6757 5363
rect -6683 5317 -6637 5363
rect -6563 5317 -6517 5363
rect -6443 5317 -6397 5363
rect -6323 5317 -6277 5363
rect -6203 5317 -6157 5363
rect -6083 5317 -6037 5363
<< polysilicon >>
rect -6960 6120 -6840 6180
rect -6720 6120 -6600 6180
rect -6480 6120 -6360 6180
rect -6240 6120 -6120 6180
rect -6960 5640 -6840 5760
rect -6720 5640 -6600 5760
rect -6480 5640 -6360 5760
rect -6240 5640 -6120 5760
rect -6960 5603 -6120 5640
rect -6960 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6563 5603
rect -6517 5557 -6443 5603
rect -6397 5557 -6323 5603
rect -6277 5557 -6203 5603
rect -6157 5557 -6120 5603
rect -6960 5520 -6120 5557
rect -6960 4500 -6840 4560
rect -6720 4500 -6600 4560
rect -6480 4500 -6360 4560
rect -6240 4500 -6120 4560
rect -6960 4080 -6840 4200
rect -6720 4080 -6600 4200
rect -6960 4043 -6600 4080
rect -6960 3997 -6923 4043
rect -6877 3997 -6803 4043
rect -6757 3997 -6683 4043
rect -6637 3997 -6600 4043
rect -6960 3960 -6600 3997
rect -6480 4080 -6360 4200
rect -6240 4080 -6120 4200
rect -6480 4043 -6120 4080
rect -6480 3997 -6443 4043
rect -6397 3997 -6323 4043
rect -6277 3997 -6203 4043
rect -6157 3997 -6120 4043
rect -6480 3960 -6120 3997
rect -6960 -517 -6600 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6803 -517
rect -6757 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -600 -6600 -563
rect -6960 -720 -6840 -600
rect -6720 -720 -6600 -600
rect -6480 -517 -6120 -480
rect -6480 -563 -6443 -517
rect -6397 -563 -6323 -517
rect -6277 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -600 -6120 -563
rect -6480 -720 -6360 -600
rect -6240 -720 -6120 -600
rect -6960 -1140 -6840 -1080
rect -6720 -1140 -6600 -1080
rect -6480 -1140 -6360 -1080
rect -6240 -1140 -6120 -1080
<< polycontact >>
rect -6923 5557 -6877 5603
rect -6803 5557 -6757 5603
rect -6683 5557 -6637 5603
rect -6563 5557 -6517 5603
rect -6443 5557 -6397 5603
rect -6323 5557 -6277 5603
rect -6203 5557 -6157 5603
rect -6923 3997 -6877 4043
rect -6803 3997 -6757 4043
rect -6683 3997 -6637 4043
rect -6443 3997 -6397 4043
rect -6323 3997 -6277 4043
rect -6203 3997 -6157 4043
rect -6923 -563 -6877 -517
rect -6803 -563 -6757 -517
rect -6683 -563 -6637 -517
rect -6443 -563 -6397 -517
rect -6323 -563 -6277 -517
rect -6203 -563 -6157 -517
<< metal1 >>
rect -7200 6563 -5880 6600
rect -7200 6517 -7163 6563
rect -7117 6517 -7043 6563
rect -6997 6517 -6923 6563
rect -6877 6517 -6803 6563
rect -6757 6517 -6683 6563
rect -6637 6517 -6563 6563
rect -6517 6517 -6443 6563
rect -6397 6517 -6323 6563
rect -6277 6517 -6203 6563
rect -6157 6517 -6083 6563
rect -6037 6517 -5963 6563
rect -5917 6517 -5880 6563
rect -7200 6480 -5880 6517
rect -7200 6326 -5880 6360
rect -7200 6274 -7046 6326
rect -6994 6323 -6566 6326
rect -6514 6323 -6086 6326
rect -6994 6277 -6923 6323
rect -6877 6277 -6803 6323
rect -6757 6277 -6683 6323
rect -6637 6277 -6566 6323
rect -6514 6277 -6443 6323
rect -6397 6277 -6323 6323
rect -6277 6277 -6203 6323
rect -6157 6277 -6086 6323
rect -6994 6274 -6566 6277
rect -6514 6274 -6086 6277
rect -6034 6274 -5880 6326
rect -7200 6240 -5880 6274
rect -7080 6086 -6960 6120
rect -7080 6034 -7046 6086
rect -6994 6034 -6960 6086
rect -7080 5966 -6960 6034
rect -7080 5914 -7046 5966
rect -6994 5914 -6960 5966
rect -7080 5846 -6960 5914
rect -7080 5794 -7046 5846
rect -6994 5794 -6960 5846
rect -7080 5760 -6960 5794
rect -6840 6086 -6720 6120
rect -6840 6034 -6806 6086
rect -6754 6034 -6720 6086
rect -6840 5966 -6720 6034
rect -6840 5914 -6806 5966
rect -6754 5914 -6720 5966
rect -6840 5846 -6720 5914
rect -6840 5794 -6806 5846
rect -6754 5794 -6720 5846
rect -6840 5760 -6720 5794
rect -6600 6086 -6480 6120
rect -6600 6034 -6566 6086
rect -6514 6034 -6480 6086
rect -6600 5966 -6480 6034
rect -6600 5914 -6566 5966
rect -6514 5914 -6480 5966
rect -6600 5846 -6480 5914
rect -6600 5794 -6566 5846
rect -6514 5794 -6480 5846
rect -6600 5760 -6480 5794
rect -6360 6086 -6240 6120
rect -6360 6034 -6326 6086
rect -6274 6034 -6240 6086
rect -6360 5966 -6240 6034
rect -6360 5914 -6326 5966
rect -6274 5914 -6240 5966
rect -6360 5846 -6240 5914
rect -6360 5794 -6326 5846
rect -6274 5794 -6240 5846
rect -6360 5760 -6240 5794
rect -6120 6086 -6000 6120
rect -6120 6034 -6086 6086
rect -6034 6034 -6000 6086
rect -6120 5966 -6000 6034
rect -6120 5914 -6086 5966
rect -6034 5914 -6000 5966
rect -6120 5846 -6000 5914
rect -6120 5794 -6086 5846
rect -6034 5794 -6000 5846
rect -6120 5760 -6000 5794
rect -6960 5606 -6120 5640
rect -6960 5603 -6566 5606
rect -6514 5603 -6120 5606
rect -6960 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6566 5603
rect -6514 5557 -6443 5603
rect -6397 5557 -6323 5603
rect -6277 5557 -6203 5603
rect -6157 5557 -6120 5603
rect -6960 5554 -6566 5557
rect -6514 5554 -6120 5557
rect -6960 5520 -6120 5554
rect -7200 5363 -5880 5400
rect -7200 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6683 5363
rect -6637 5317 -6563 5363
rect -6517 5317 -6443 5363
rect -6397 5317 -6323 5363
rect -6277 5317 -6203 5363
rect -6157 5317 -6083 5363
rect -6037 5317 -5880 5363
rect -7200 5280 -5880 5317
rect -7200 5123 -5880 5160
rect -7200 5077 -7163 5123
rect -7117 5077 -7043 5123
rect -6997 5077 -6923 5123
rect -6877 5077 -6803 5123
rect -6757 5077 -6683 5123
rect -6637 5077 -6563 5123
rect -6517 5077 -6443 5123
rect -6397 5077 -6323 5123
rect -6277 5077 -6203 5123
rect -6157 5077 -6083 5123
rect -6037 5077 -5963 5123
rect -5917 5077 -5880 5123
rect -7200 5040 -5880 5077
rect -7200 4883 -5880 4920
rect -7200 4837 -7043 4883
rect -6997 4837 -6923 4883
rect -6877 4837 -6803 4883
rect -6757 4837 -6683 4883
rect -6637 4837 -6563 4883
rect -6517 4837 -6443 4883
rect -6397 4837 -6323 4883
rect -6277 4837 -6203 4883
rect -6157 4837 -6083 4883
rect -6037 4837 -5880 4883
rect -7200 4800 -5880 4837
rect -7080 4646 -6000 4680
rect -7080 4594 -7046 4646
rect -6994 4594 -6566 4646
rect -6514 4594 -6086 4646
rect -6034 4594 -6000 4646
rect -7080 4560 -6000 4594
rect -7080 4526 -6960 4560
rect -7080 4474 -7046 4526
rect -6994 4474 -6960 4526
rect -6600 4526 -6480 4560
rect -7080 4406 -6960 4474
rect -7080 4354 -7046 4406
rect -6994 4354 -6960 4406
rect -7080 4286 -6960 4354
rect -7080 4234 -7046 4286
rect -6994 4234 -6960 4286
rect -7080 4200 -6960 4234
rect -6840 4406 -6720 4500
rect -6840 4354 -6806 4406
rect -6754 4354 -6720 4406
rect -6840 4286 -6720 4354
rect -6840 4234 -6806 4286
rect -6754 4234 -6720 4286
rect -6840 4200 -6720 4234
rect -6600 4474 -6566 4526
rect -6514 4474 -6480 4526
rect -6120 4526 -6000 4560
rect -6600 4403 -6480 4474
rect -6600 4357 -6563 4403
rect -6517 4357 -6480 4403
rect -6600 4283 -6480 4357
rect -6600 4237 -6563 4283
rect -6517 4237 -6480 4283
rect -6600 4200 -6480 4237
rect -6360 4406 -6240 4500
rect -6360 4354 -6326 4406
rect -6274 4354 -6240 4406
rect -6360 4286 -6240 4354
rect -6360 4234 -6326 4286
rect -6274 4234 -6240 4286
rect -6360 4200 -6240 4234
rect -6120 4474 -6086 4526
rect -6034 4474 -6000 4526
rect -6120 4406 -6000 4474
rect -6120 4354 -6086 4406
rect -6034 4354 -6000 4406
rect -6120 4286 -6000 4354
rect -6120 4234 -6086 4286
rect -6034 4234 -6000 4286
rect -6120 4200 -6000 4234
rect -6960 4046 -6600 4080
rect -6960 4043 -6806 4046
rect -6754 4043 -6600 4046
rect -6960 3997 -6923 4043
rect -6877 3997 -6806 4043
rect -6754 3997 -6683 4043
rect -6637 3997 -6600 4043
rect -6960 3994 -6806 3997
rect -6754 3994 -6600 3997
rect -6960 3960 -6600 3994
rect -6480 4046 -6120 4080
rect -6480 4043 -6326 4046
rect -6274 4043 -6120 4046
rect -6480 3997 -6443 4043
rect -6397 3997 -6326 4043
rect -6274 3997 -6203 4043
rect -6157 3997 -6120 4043
rect -6480 3994 -6326 3997
rect -6274 3994 -6120 3997
rect -6480 3960 -6120 3994
rect -7200 3806 -5880 3840
rect -7200 3754 -7046 3806
rect -6994 3803 -6086 3806
rect -6994 3757 -6923 3803
rect -6877 3757 -6803 3803
rect -6757 3757 -6683 3803
rect -6637 3757 -6563 3803
rect -6517 3757 -6443 3803
rect -6397 3757 -6323 3803
rect -6277 3757 -6203 3803
rect -6157 3757 -6086 3803
rect -6994 3754 -6086 3757
rect -6034 3754 -5880 3806
rect -7200 3720 -5880 3754
rect -7200 3566 -5880 3600
rect -7200 3563 -7046 3566
rect -6994 3563 -6086 3566
rect -6034 3563 -5880 3566
rect -7200 3517 -7163 3563
rect -7117 3517 -7046 3563
rect -6994 3517 -6923 3563
rect -6877 3517 -6803 3563
rect -6757 3517 -6683 3563
rect -6637 3517 -6563 3563
rect -6517 3517 -6443 3563
rect -6397 3517 -6323 3563
rect -6277 3517 -6203 3563
rect -6157 3517 -6086 3563
rect -6034 3517 -5963 3563
rect -5917 3517 -5880 3563
rect -7200 3514 -7046 3517
rect -6994 3514 -6086 3517
rect -6034 3514 -5880 3517
rect -7200 3480 -5880 3514
rect -7200 2606 -5880 2640
rect -7200 2603 -7046 2606
rect -6994 2603 -6086 2606
rect -6034 2603 -5880 2606
rect -7200 2557 -7163 2603
rect -7117 2557 -7046 2603
rect -6994 2557 -6923 2603
rect -6877 2557 -6803 2603
rect -6757 2557 -6683 2603
rect -6637 2557 -6563 2603
rect -6517 2557 -6443 2603
rect -6397 2557 -6323 2603
rect -6277 2557 -6203 2603
rect -6157 2557 -6086 2603
rect -6034 2557 -5963 2603
rect -5917 2557 -5880 2603
rect -7200 2554 -7046 2557
rect -6994 2554 -6086 2557
rect -6034 2554 -5880 2557
rect -7200 2520 -5880 2554
rect -7200 2126 -5880 2160
rect -7200 2123 -7046 2126
rect -6994 2123 -6086 2126
rect -6034 2123 -5880 2126
rect -7200 2077 -7163 2123
rect -7117 2077 -7046 2123
rect -6994 2077 -6923 2123
rect -6877 2077 -6803 2123
rect -6757 2077 -6683 2123
rect -6637 2077 -6563 2123
rect -6517 2077 -6443 2123
rect -6397 2077 -6323 2123
rect -6277 2077 -6203 2123
rect -6157 2077 -6086 2123
rect -6034 2077 -5963 2123
rect -5917 2077 -5880 2123
rect -7200 2074 -7046 2077
rect -6994 2074 -6086 2077
rect -6034 2074 -5880 2077
rect -7200 2040 -5880 2074
rect -7200 1646 -5880 1680
rect -7200 1643 -7046 1646
rect -6994 1643 -6086 1646
rect -6034 1643 -5880 1646
rect -7200 1597 -7163 1643
rect -7117 1597 -7046 1643
rect -6994 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6563 1643
rect -6517 1597 -6443 1643
rect -6397 1597 -6323 1643
rect -6277 1597 -6203 1643
rect -6157 1597 -6086 1643
rect -6034 1597 -5963 1643
rect -5917 1597 -5880 1643
rect -7200 1594 -7046 1597
rect -6994 1594 -6086 1597
rect -6034 1594 -5880 1597
rect -7200 1560 -5880 1594
rect -7200 1166 -5880 1200
rect -7200 1163 -7046 1166
rect -6994 1163 -6086 1166
rect -6034 1163 -5880 1166
rect -7200 1117 -7163 1163
rect -7117 1117 -7046 1163
rect -6994 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6563 1163
rect -6517 1117 -6443 1163
rect -6397 1117 -6323 1163
rect -6277 1117 -6203 1163
rect -6157 1117 -6086 1163
rect -6034 1117 -5963 1163
rect -5917 1117 -5880 1163
rect -7200 1114 -7046 1117
rect -6994 1114 -6086 1117
rect -6034 1114 -5880 1117
rect -7200 1080 -5880 1114
rect -7200 686 -5880 720
rect -7200 683 -7046 686
rect -6994 683 -6086 686
rect -6034 683 -5880 686
rect -7200 637 -7163 683
rect -7117 637 -7046 683
rect -6994 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6563 683
rect -6517 637 -6443 683
rect -6397 637 -6323 683
rect -6277 637 -6203 683
rect -6157 637 -6086 683
rect -6034 637 -5963 683
rect -5917 637 -5880 683
rect -7200 634 -7046 637
rect -6994 634 -6086 637
rect -6034 634 -5880 637
rect -7200 600 -5880 634
rect -7200 -274 -5880 -240
rect -7200 -277 -7046 -274
rect -6994 -277 -6086 -274
rect -6034 -277 -5880 -274
rect -7200 -323 -7163 -277
rect -7117 -323 -7046 -277
rect -6994 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6086 -277
rect -6034 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -326 -7046 -323
rect -6994 -326 -6086 -323
rect -6034 -326 -5880 -323
rect -7200 -360 -5880 -326
rect -6960 -514 -6600 -480
rect -6960 -517 -6806 -514
rect -6754 -517 -6600 -514
rect -6960 -563 -6923 -517
rect -6877 -563 -6806 -517
rect -6754 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -566 -6806 -563
rect -6754 -566 -6600 -563
rect -6960 -600 -6600 -566
rect -6480 -514 -6120 -480
rect -6480 -517 -6326 -514
rect -6274 -517 -6120 -514
rect -6480 -563 -6443 -517
rect -6397 -563 -6326 -517
rect -6274 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -566 -6326 -563
rect -6274 -566 -6120 -563
rect -6480 -600 -6120 -566
rect -7080 -754 -6960 -720
rect -7080 -806 -7046 -754
rect -6994 -806 -6960 -754
rect -7080 -874 -6960 -806
rect -7080 -926 -7046 -874
rect -6994 -926 -6960 -874
rect -7080 -994 -6960 -926
rect -7080 -1046 -7046 -994
rect -6994 -1046 -6960 -994
rect -7080 -1080 -6960 -1046
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -754 -6480 -720
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -754 -6000 -720
rect -6120 -806 -6086 -754
rect -6034 -806 -6000 -754
rect -6120 -874 -6000 -806
rect -6120 -926 -6086 -874
rect -6034 -926 -6000 -874
rect -6120 -994 -6000 -926
rect -6120 -1046 -6086 -994
rect -6034 -1046 -6000 -994
rect -6120 -1080 -6000 -1046
rect -7200 -1234 -5880 -1200
rect -7200 -1237 -7046 -1234
rect -6994 -1237 -6086 -1234
rect -6034 -1237 -5880 -1234
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7046 -1237
rect -6994 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6086 -1237
rect -6034 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1286 -7046 -1283
rect -6994 -1286 -6086 -1283
rect -6034 -1286 -5880 -1283
rect -7200 -1320 -5880 -1286
<< via1 >>
rect -7046 6323 -6994 6326
rect -6566 6323 -6514 6326
rect -6086 6323 -6034 6326
rect -7046 6277 -7043 6323
rect -7043 6277 -6997 6323
rect -6997 6277 -6994 6323
rect -6566 6277 -6563 6323
rect -6563 6277 -6517 6323
rect -6517 6277 -6514 6323
rect -6086 6277 -6083 6323
rect -6083 6277 -6037 6323
rect -6037 6277 -6034 6323
rect -7046 6274 -6994 6277
rect -6566 6274 -6514 6277
rect -6086 6274 -6034 6277
rect -7046 6083 -6994 6086
rect -7046 6037 -7043 6083
rect -7043 6037 -6997 6083
rect -6997 6037 -6994 6083
rect -7046 6034 -6994 6037
rect -7046 5963 -6994 5966
rect -7046 5917 -7043 5963
rect -7043 5917 -6997 5963
rect -6997 5917 -6994 5963
rect -7046 5914 -6994 5917
rect -7046 5843 -6994 5846
rect -7046 5797 -7043 5843
rect -7043 5797 -6997 5843
rect -6997 5797 -6994 5843
rect -7046 5794 -6994 5797
rect -6806 6083 -6754 6086
rect -6806 6037 -6803 6083
rect -6803 6037 -6757 6083
rect -6757 6037 -6754 6083
rect -6806 6034 -6754 6037
rect -6806 5963 -6754 5966
rect -6806 5917 -6803 5963
rect -6803 5917 -6757 5963
rect -6757 5917 -6754 5963
rect -6806 5914 -6754 5917
rect -6806 5843 -6754 5846
rect -6806 5797 -6803 5843
rect -6803 5797 -6757 5843
rect -6757 5797 -6754 5843
rect -6806 5794 -6754 5797
rect -6566 6083 -6514 6086
rect -6566 6037 -6563 6083
rect -6563 6037 -6517 6083
rect -6517 6037 -6514 6083
rect -6566 6034 -6514 6037
rect -6566 5963 -6514 5966
rect -6566 5917 -6563 5963
rect -6563 5917 -6517 5963
rect -6517 5917 -6514 5963
rect -6566 5914 -6514 5917
rect -6566 5843 -6514 5846
rect -6566 5797 -6563 5843
rect -6563 5797 -6517 5843
rect -6517 5797 -6514 5843
rect -6566 5794 -6514 5797
rect -6326 6083 -6274 6086
rect -6326 6037 -6323 6083
rect -6323 6037 -6277 6083
rect -6277 6037 -6274 6083
rect -6326 6034 -6274 6037
rect -6326 5963 -6274 5966
rect -6326 5917 -6323 5963
rect -6323 5917 -6277 5963
rect -6277 5917 -6274 5963
rect -6326 5914 -6274 5917
rect -6326 5843 -6274 5846
rect -6326 5797 -6323 5843
rect -6323 5797 -6277 5843
rect -6277 5797 -6274 5843
rect -6326 5794 -6274 5797
rect -6086 6083 -6034 6086
rect -6086 6037 -6083 6083
rect -6083 6037 -6037 6083
rect -6037 6037 -6034 6083
rect -6086 6034 -6034 6037
rect -6086 5963 -6034 5966
rect -6086 5917 -6083 5963
rect -6083 5917 -6037 5963
rect -6037 5917 -6034 5963
rect -6086 5914 -6034 5917
rect -6086 5843 -6034 5846
rect -6086 5797 -6083 5843
rect -6083 5797 -6037 5843
rect -6037 5797 -6034 5843
rect -6086 5794 -6034 5797
rect -6566 5603 -6514 5606
rect -6566 5557 -6563 5603
rect -6563 5557 -6517 5603
rect -6517 5557 -6514 5603
rect -6566 5554 -6514 5557
rect -7046 4594 -6994 4646
rect -6566 4594 -6514 4646
rect -6086 4594 -6034 4646
rect -7046 4474 -6994 4526
rect -7046 4403 -6994 4406
rect -7046 4357 -7043 4403
rect -7043 4357 -6997 4403
rect -6997 4357 -6994 4403
rect -7046 4354 -6994 4357
rect -7046 4283 -6994 4286
rect -7046 4237 -7043 4283
rect -7043 4237 -6997 4283
rect -6997 4237 -6994 4283
rect -7046 4234 -6994 4237
rect -6806 4403 -6754 4406
rect -6806 4357 -6803 4403
rect -6803 4357 -6757 4403
rect -6757 4357 -6754 4403
rect -6806 4354 -6754 4357
rect -6806 4283 -6754 4286
rect -6806 4237 -6803 4283
rect -6803 4237 -6757 4283
rect -6757 4237 -6754 4283
rect -6806 4234 -6754 4237
rect -6566 4474 -6514 4526
rect -6326 4403 -6274 4406
rect -6326 4357 -6323 4403
rect -6323 4357 -6277 4403
rect -6277 4357 -6274 4403
rect -6326 4354 -6274 4357
rect -6326 4283 -6274 4286
rect -6326 4237 -6323 4283
rect -6323 4237 -6277 4283
rect -6277 4237 -6274 4283
rect -6326 4234 -6274 4237
rect -6086 4474 -6034 4526
rect -6086 4403 -6034 4406
rect -6086 4357 -6083 4403
rect -6083 4357 -6037 4403
rect -6037 4357 -6034 4403
rect -6086 4354 -6034 4357
rect -6086 4283 -6034 4286
rect -6086 4237 -6083 4283
rect -6083 4237 -6037 4283
rect -6037 4237 -6034 4283
rect -6086 4234 -6034 4237
rect -6806 4043 -6754 4046
rect -6806 3997 -6803 4043
rect -6803 3997 -6757 4043
rect -6757 3997 -6754 4043
rect -6806 3994 -6754 3997
rect -6326 4043 -6274 4046
rect -6326 3997 -6323 4043
rect -6323 3997 -6277 4043
rect -6277 3997 -6274 4043
rect -6326 3994 -6274 3997
rect -7046 3803 -6994 3806
rect -6086 3803 -6034 3806
rect -7046 3757 -7043 3803
rect -7043 3757 -6997 3803
rect -6997 3757 -6994 3803
rect -6086 3757 -6083 3803
rect -6083 3757 -6037 3803
rect -6037 3757 -6034 3803
rect -7046 3754 -6994 3757
rect -6086 3754 -6034 3757
rect -7046 3563 -6994 3566
rect -6086 3563 -6034 3566
rect -7046 3517 -7043 3563
rect -7043 3517 -6997 3563
rect -6997 3517 -6994 3563
rect -6086 3517 -6083 3563
rect -6083 3517 -6037 3563
rect -6037 3517 -6034 3563
rect -7046 3514 -6994 3517
rect -6086 3514 -6034 3517
rect -7046 2603 -6994 2606
rect -6086 2603 -6034 2606
rect -7046 2557 -7043 2603
rect -7043 2557 -6997 2603
rect -6997 2557 -6994 2603
rect -6086 2557 -6083 2603
rect -6083 2557 -6037 2603
rect -6037 2557 -6034 2603
rect -7046 2554 -6994 2557
rect -6086 2554 -6034 2557
rect -7046 2123 -6994 2126
rect -6086 2123 -6034 2126
rect -7046 2077 -7043 2123
rect -7043 2077 -6997 2123
rect -6997 2077 -6994 2123
rect -6086 2077 -6083 2123
rect -6083 2077 -6037 2123
rect -6037 2077 -6034 2123
rect -7046 2074 -6994 2077
rect -6086 2074 -6034 2077
rect -7046 1643 -6994 1646
rect -6086 1643 -6034 1646
rect -7046 1597 -7043 1643
rect -7043 1597 -6997 1643
rect -6997 1597 -6994 1643
rect -6086 1597 -6083 1643
rect -6083 1597 -6037 1643
rect -6037 1597 -6034 1643
rect -7046 1594 -6994 1597
rect -6086 1594 -6034 1597
rect -7046 1163 -6994 1166
rect -6086 1163 -6034 1166
rect -7046 1117 -7043 1163
rect -7043 1117 -6997 1163
rect -6997 1117 -6994 1163
rect -6086 1117 -6083 1163
rect -6083 1117 -6037 1163
rect -6037 1117 -6034 1163
rect -7046 1114 -6994 1117
rect -6086 1114 -6034 1117
rect -7046 683 -6994 686
rect -6086 683 -6034 686
rect -7046 637 -7043 683
rect -7043 637 -6997 683
rect -6997 637 -6994 683
rect -6086 637 -6083 683
rect -6083 637 -6037 683
rect -6037 637 -6034 683
rect -7046 634 -6994 637
rect -6086 634 -6034 637
rect -7046 -277 -6994 -274
rect -6086 -277 -6034 -274
rect -7046 -323 -7043 -277
rect -7043 -323 -6997 -277
rect -6997 -323 -6994 -277
rect -6086 -323 -6083 -277
rect -6083 -323 -6037 -277
rect -6037 -323 -6034 -277
rect -7046 -326 -6994 -323
rect -6086 -326 -6034 -323
rect -6806 -517 -6754 -514
rect -6806 -563 -6803 -517
rect -6803 -563 -6757 -517
rect -6757 -563 -6754 -517
rect -6806 -566 -6754 -563
rect -6326 -517 -6274 -514
rect -6326 -563 -6323 -517
rect -6323 -563 -6277 -517
rect -6277 -563 -6274 -517
rect -6326 -566 -6274 -563
rect -7046 -757 -6994 -754
rect -7046 -803 -7043 -757
rect -7043 -803 -6997 -757
rect -6997 -803 -6994 -757
rect -7046 -806 -6994 -803
rect -7046 -877 -6994 -874
rect -7046 -923 -7043 -877
rect -7043 -923 -6997 -877
rect -6997 -923 -6994 -877
rect -7046 -926 -6994 -923
rect -7046 -997 -6994 -994
rect -7046 -1043 -7043 -997
rect -7043 -1043 -6997 -997
rect -6997 -1043 -6994 -997
rect -7046 -1046 -6994 -1043
rect -6566 -757 -6514 -754
rect -6566 -803 -6563 -757
rect -6563 -803 -6517 -757
rect -6517 -803 -6514 -757
rect -6566 -806 -6514 -803
rect -6566 -877 -6514 -874
rect -6566 -923 -6563 -877
rect -6563 -923 -6517 -877
rect -6517 -923 -6514 -877
rect -6566 -926 -6514 -923
rect -6566 -997 -6514 -994
rect -6566 -1043 -6563 -997
rect -6563 -1043 -6517 -997
rect -6517 -1043 -6514 -997
rect -6566 -1046 -6514 -1043
rect -6086 -757 -6034 -754
rect -6086 -803 -6083 -757
rect -6083 -803 -6037 -757
rect -6037 -803 -6034 -757
rect -6086 -806 -6034 -803
rect -6086 -877 -6034 -874
rect -6086 -923 -6083 -877
rect -6083 -923 -6037 -877
rect -6037 -923 -6034 -877
rect -6086 -926 -6034 -923
rect -6086 -997 -6034 -994
rect -6086 -1043 -6083 -997
rect -6083 -1043 -6037 -997
rect -6037 -1043 -6034 -997
rect -6086 -1046 -6034 -1043
rect -7046 -1237 -6994 -1234
rect -6086 -1237 -6034 -1234
rect -7046 -1283 -7043 -1237
rect -7043 -1283 -6997 -1237
rect -6997 -1283 -6994 -1237
rect -6086 -1283 -6083 -1237
rect -6083 -1283 -6037 -1237
rect -6037 -1283 -6034 -1237
rect -7046 -1286 -6994 -1283
rect -6086 -1286 -6034 -1283
<< metal2 >>
rect -7080 6328 -6960 6360
rect -7080 6272 -7048 6328
rect -6992 6272 -6960 6328
rect -7080 6088 -6960 6272
rect -6600 6328 -6480 6360
rect -6600 6272 -6568 6328
rect -6512 6272 -6480 6328
rect -7080 6032 -7048 6088
rect -6992 6032 -6960 6088
rect -7080 5968 -6960 6032
rect -7080 5912 -7048 5968
rect -6992 5912 -6960 5968
rect -7080 5848 -6960 5912
rect -7080 5792 -7048 5848
rect -6992 5792 -6960 5848
rect -7080 5760 -6960 5792
rect -6840 6086 -6720 6120
rect -6840 6034 -6806 6086
rect -6754 6034 -6720 6086
rect -6840 5966 -6720 6034
rect -6840 5914 -6806 5966
rect -6754 5914 -6720 5966
rect -6840 5846 -6720 5914
rect -6840 5794 -6806 5846
rect -6754 5794 -6720 5846
rect -6840 5368 -6720 5794
rect -6600 6088 -6480 6272
rect -6120 6328 -6000 6360
rect -6120 6272 -6088 6328
rect -6032 6272 -6000 6328
rect -6600 6032 -6568 6088
rect -6512 6032 -6480 6088
rect -6600 5968 -6480 6032
rect -6600 5912 -6568 5968
rect -6512 5912 -6480 5968
rect -6600 5848 -6480 5912
rect -6600 5792 -6568 5848
rect -6512 5792 -6480 5848
rect -6600 5760 -6480 5792
rect -6360 6086 -6240 6120
rect -6360 6034 -6326 6086
rect -6274 6034 -6240 6086
rect -6360 5966 -6240 6034
rect -6360 5914 -6326 5966
rect -6274 5914 -6240 5966
rect -6360 5846 -6240 5914
rect -6360 5794 -6326 5846
rect -6274 5794 -6240 5846
rect -6600 5608 -6480 5640
rect -6600 5552 -6568 5608
rect -6512 5552 -6480 5608
rect -6600 5520 -6480 5552
rect -6840 5312 -6808 5368
rect -6752 5312 -6720 5368
rect -7080 4888 -6960 4920
rect -7080 4832 -7048 4888
rect -6992 4832 -6960 4888
rect -7080 4646 -6960 4832
rect -6840 4888 -6720 5312
rect -6360 5368 -6240 5794
rect -6120 6088 -6000 6272
rect -6120 6032 -6088 6088
rect -6032 6032 -6000 6088
rect -6120 5968 -6000 6032
rect -6120 5912 -6088 5968
rect -6032 5912 -6000 5968
rect -6120 5848 -6000 5912
rect -6120 5792 -6088 5848
rect -6032 5792 -6000 5848
rect -6120 5760 -6000 5792
rect -6360 5312 -6328 5368
rect -6272 5312 -6240 5368
rect -6840 4832 -6808 4888
rect -6752 4832 -6720 4888
rect -6840 4800 -6720 4832
rect -6600 4888 -6480 4920
rect -6600 4832 -6568 4888
rect -6512 4832 -6480 4888
rect -7080 4594 -7046 4646
rect -6994 4594 -6960 4646
rect -7080 4526 -6960 4594
rect -7080 4474 -7046 4526
rect -6994 4474 -6960 4526
rect -6600 4646 -6480 4832
rect -6360 4888 -6240 5312
rect -6360 4832 -6328 4888
rect -6272 4832 -6240 4888
rect -6360 4800 -6240 4832
rect -6120 4888 -6000 4920
rect -6120 4832 -6088 4888
rect -6032 4832 -6000 4888
rect -6600 4594 -6566 4646
rect -6514 4594 -6480 4646
rect -6600 4526 -6480 4594
rect -7080 4406 -6960 4474
rect -7080 4354 -7046 4406
rect -6994 4354 -6960 4406
rect -7080 4286 -6960 4354
rect -7080 4234 -7046 4286
rect -6994 4234 -6960 4286
rect -7080 4200 -6960 4234
rect -6840 4406 -6720 4500
rect -6600 4474 -6566 4526
rect -6514 4474 -6480 4526
rect -6120 4646 -6000 4832
rect -6120 4594 -6086 4646
rect -6034 4594 -6000 4646
rect -6120 4526 -6000 4594
rect -6600 4440 -6480 4474
rect -6840 4354 -6806 4406
rect -6754 4354 -6720 4406
rect -6840 4320 -6720 4354
rect -6360 4406 -6240 4500
rect -6360 4354 -6326 4406
rect -6274 4354 -6240 4406
rect -6360 4320 -6240 4354
rect -6840 4286 -6240 4320
rect -6840 4234 -6806 4286
rect -6754 4234 -6326 4286
rect -6274 4234 -6240 4286
rect -6840 4200 -6240 4234
rect -6120 4474 -6086 4526
rect -6034 4474 -6000 4526
rect -6120 4406 -6000 4474
rect -6120 4354 -6086 4406
rect -6034 4354 -6000 4406
rect -6120 4286 -6000 4354
rect -6120 4234 -6086 4286
rect -6034 4234 -6000 4286
rect -6120 4200 -6000 4234
rect -6840 4048 -6720 4080
rect -6840 3992 -6808 4048
rect -6752 3992 -6720 4048
rect -6840 3960 -6720 3992
rect -7080 3808 -6960 3840
rect -7080 3752 -7048 3808
rect -6992 3752 -6960 3808
rect -7080 3720 -6960 3752
rect -7080 3568 -6960 3600
rect -7080 3512 -7048 3568
rect -6992 3512 -6960 3568
rect -7080 2608 -6960 3512
rect -7080 2552 -7048 2608
rect -6992 2552 -6960 2608
rect -7080 2128 -6960 2552
rect -7080 2072 -7048 2128
rect -6992 2072 -6960 2128
rect -7080 1648 -6960 2072
rect -7080 1592 -7048 1648
rect -6992 1592 -6960 1648
rect -7080 1168 -6960 1592
rect -7080 1112 -7048 1168
rect -6992 1112 -6960 1168
rect -7080 688 -6960 1112
rect -7080 632 -7048 688
rect -6992 632 -6960 688
rect -7080 -272 -6960 632
rect -7080 -328 -7048 -272
rect -6992 -328 -6960 -272
rect -7080 -752 -6960 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -7080 -808 -7048 -752
rect -6992 -808 -6960 -752
rect -7080 -872 -6960 -808
rect -7080 -928 -7048 -872
rect -6992 -928 -6960 -872
rect -7080 -992 -6960 -928
rect -7080 -1048 -7048 -992
rect -6992 -1048 -6960 -992
rect -7080 -1232 -6960 -1048
rect -6600 -754 -6480 4200
rect -6360 4048 -6240 4080
rect -6360 3992 -6328 4048
rect -6272 3992 -6240 4048
rect -6360 3960 -6240 3992
rect -6120 3808 -6000 3840
rect -6120 3752 -6088 3808
rect -6032 3752 -6000 3808
rect -6120 3720 -6000 3752
rect -6120 3568 -6000 3600
rect -6120 3512 -6088 3568
rect -6032 3512 -6000 3568
rect -6120 2608 -6000 3512
rect -6120 2552 -6088 2608
rect -6032 2552 -6000 2608
rect -6120 2128 -6000 2552
rect -6120 2072 -6088 2128
rect -6032 2072 -6000 2128
rect -6120 1648 -6000 2072
rect -6120 1592 -6088 1648
rect -6032 1592 -6000 1648
rect -6120 1168 -6000 1592
rect -6120 1112 -6088 1168
rect -6032 1112 -6000 1168
rect -6120 688 -6000 1112
rect -6120 632 -6088 688
rect -6032 632 -6000 688
rect -6120 -272 -6000 632
rect -6120 -328 -6088 -272
rect -6032 -328 -6000 -272
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6120 -752 -6000 -328
rect -6120 -808 -6088 -752
rect -6032 -808 -6000 -752
rect -6120 -872 -6000 -808
rect -6120 -928 -6088 -872
rect -6032 -928 -6000 -872
rect -6120 -992 -6000 -928
rect -6120 -1048 -6088 -992
rect -6032 -1048 -6000 -992
rect -7080 -1288 -7048 -1232
rect -6992 -1288 -6960 -1232
rect -7080 -1320 -6960 -1288
rect -6120 -1232 -6000 -1048
rect -6120 -1288 -6088 -1232
rect -6032 -1288 -6000 -1232
rect -6120 -1320 -6000 -1288
<< via2 >>
rect -7048 6326 -6992 6328
rect -7048 6274 -7046 6326
rect -7046 6274 -6994 6326
rect -6994 6274 -6992 6326
rect -7048 6272 -6992 6274
rect -6568 6326 -6512 6328
rect -6568 6274 -6566 6326
rect -6566 6274 -6514 6326
rect -6514 6274 -6512 6326
rect -6568 6272 -6512 6274
rect -7048 6086 -6992 6088
rect -7048 6034 -7046 6086
rect -7046 6034 -6994 6086
rect -6994 6034 -6992 6086
rect -7048 6032 -6992 6034
rect -7048 5966 -6992 5968
rect -7048 5914 -7046 5966
rect -7046 5914 -6994 5966
rect -6994 5914 -6992 5966
rect -7048 5912 -6992 5914
rect -7048 5846 -6992 5848
rect -7048 5794 -7046 5846
rect -7046 5794 -6994 5846
rect -6994 5794 -6992 5846
rect -7048 5792 -6992 5794
rect -6088 6326 -6032 6328
rect -6088 6274 -6086 6326
rect -6086 6274 -6034 6326
rect -6034 6274 -6032 6326
rect -6088 6272 -6032 6274
rect -6568 6086 -6512 6088
rect -6568 6034 -6566 6086
rect -6566 6034 -6514 6086
rect -6514 6034 -6512 6086
rect -6568 6032 -6512 6034
rect -6568 5966 -6512 5968
rect -6568 5914 -6566 5966
rect -6566 5914 -6514 5966
rect -6514 5914 -6512 5966
rect -6568 5912 -6512 5914
rect -6568 5846 -6512 5848
rect -6568 5794 -6566 5846
rect -6566 5794 -6514 5846
rect -6514 5794 -6512 5846
rect -6568 5792 -6512 5794
rect -6568 5606 -6512 5608
rect -6568 5554 -6566 5606
rect -6566 5554 -6514 5606
rect -6514 5554 -6512 5606
rect -6568 5552 -6512 5554
rect -6808 5312 -6752 5368
rect -7048 4832 -6992 4888
rect -6088 6086 -6032 6088
rect -6088 6034 -6086 6086
rect -6086 6034 -6034 6086
rect -6034 6034 -6032 6086
rect -6088 6032 -6032 6034
rect -6088 5966 -6032 5968
rect -6088 5914 -6086 5966
rect -6086 5914 -6034 5966
rect -6034 5914 -6032 5966
rect -6088 5912 -6032 5914
rect -6088 5846 -6032 5848
rect -6088 5794 -6086 5846
rect -6086 5794 -6034 5846
rect -6034 5794 -6032 5846
rect -6088 5792 -6032 5794
rect -6328 5312 -6272 5368
rect -6808 4832 -6752 4888
rect -6568 4832 -6512 4888
rect -6328 4832 -6272 4888
rect -6088 4832 -6032 4888
rect -6808 4046 -6752 4048
rect -6808 3994 -6806 4046
rect -6806 3994 -6754 4046
rect -6754 3994 -6752 4046
rect -6808 3992 -6752 3994
rect -7048 3806 -6992 3808
rect -7048 3754 -7046 3806
rect -7046 3754 -6994 3806
rect -6994 3754 -6992 3806
rect -7048 3752 -6992 3754
rect -7048 3566 -6992 3568
rect -7048 3514 -7046 3566
rect -7046 3514 -6994 3566
rect -6994 3514 -6992 3566
rect -7048 3512 -6992 3514
rect -7048 2606 -6992 2608
rect -7048 2554 -7046 2606
rect -7046 2554 -6994 2606
rect -6994 2554 -6992 2606
rect -7048 2552 -6992 2554
rect -7048 2126 -6992 2128
rect -7048 2074 -7046 2126
rect -7046 2074 -6994 2126
rect -6994 2074 -6992 2126
rect -7048 2072 -6992 2074
rect -7048 1646 -6992 1648
rect -7048 1594 -7046 1646
rect -7046 1594 -6994 1646
rect -6994 1594 -6992 1646
rect -7048 1592 -6992 1594
rect -7048 1166 -6992 1168
rect -7048 1114 -7046 1166
rect -7046 1114 -6994 1166
rect -6994 1114 -6992 1166
rect -7048 1112 -6992 1114
rect -7048 686 -6992 688
rect -7048 634 -7046 686
rect -7046 634 -6994 686
rect -6994 634 -6992 686
rect -7048 632 -6992 634
rect -7048 -274 -6992 -272
rect -7048 -326 -7046 -274
rect -7046 -326 -6994 -274
rect -6994 -326 -6992 -274
rect -7048 -328 -6992 -326
rect -6808 -514 -6752 -512
rect -6808 -566 -6806 -514
rect -6806 -566 -6754 -514
rect -6754 -566 -6752 -514
rect -6808 -568 -6752 -566
rect -7048 -754 -6992 -752
rect -7048 -806 -7046 -754
rect -7046 -806 -6994 -754
rect -6994 -806 -6992 -754
rect -7048 -808 -6992 -806
rect -7048 -874 -6992 -872
rect -7048 -926 -7046 -874
rect -7046 -926 -6994 -874
rect -6994 -926 -6992 -874
rect -7048 -928 -6992 -926
rect -7048 -994 -6992 -992
rect -7048 -1046 -7046 -994
rect -7046 -1046 -6994 -994
rect -6994 -1046 -6992 -994
rect -7048 -1048 -6992 -1046
rect -6328 4046 -6272 4048
rect -6328 3994 -6326 4046
rect -6326 3994 -6274 4046
rect -6274 3994 -6272 4046
rect -6328 3992 -6272 3994
rect -6088 3806 -6032 3808
rect -6088 3754 -6086 3806
rect -6086 3754 -6034 3806
rect -6034 3754 -6032 3806
rect -6088 3752 -6032 3754
rect -6088 3566 -6032 3568
rect -6088 3514 -6086 3566
rect -6086 3514 -6034 3566
rect -6034 3514 -6032 3566
rect -6088 3512 -6032 3514
rect -6088 2606 -6032 2608
rect -6088 2554 -6086 2606
rect -6086 2554 -6034 2606
rect -6034 2554 -6032 2606
rect -6088 2552 -6032 2554
rect -6088 2126 -6032 2128
rect -6088 2074 -6086 2126
rect -6086 2074 -6034 2126
rect -6034 2074 -6032 2126
rect -6088 2072 -6032 2074
rect -6088 1646 -6032 1648
rect -6088 1594 -6086 1646
rect -6086 1594 -6034 1646
rect -6034 1594 -6032 1646
rect -6088 1592 -6032 1594
rect -6088 1166 -6032 1168
rect -6088 1114 -6086 1166
rect -6086 1114 -6034 1166
rect -6034 1114 -6032 1166
rect -6088 1112 -6032 1114
rect -6088 686 -6032 688
rect -6088 634 -6086 686
rect -6086 634 -6034 686
rect -6034 634 -6032 686
rect -6088 632 -6032 634
rect -6088 -274 -6032 -272
rect -6088 -326 -6086 -274
rect -6086 -326 -6034 -274
rect -6034 -326 -6032 -274
rect -6088 -328 -6032 -326
rect -6328 -514 -6272 -512
rect -6328 -566 -6326 -514
rect -6326 -566 -6274 -514
rect -6274 -566 -6272 -514
rect -6328 -568 -6272 -566
rect -6088 -754 -6032 -752
rect -6088 -806 -6086 -754
rect -6086 -806 -6034 -754
rect -6034 -806 -6032 -754
rect -6088 -808 -6032 -806
rect -6088 -874 -6032 -872
rect -6088 -926 -6086 -874
rect -6086 -926 -6034 -874
rect -6034 -926 -6032 -874
rect -6088 -928 -6032 -926
rect -6088 -994 -6032 -992
rect -6088 -1046 -6086 -994
rect -6086 -1046 -6034 -994
rect -6034 -1046 -6032 -994
rect -6088 -1048 -6032 -1046
rect -7048 -1234 -6992 -1232
rect -7048 -1286 -7046 -1234
rect -7046 -1286 -6994 -1234
rect -6994 -1286 -6992 -1234
rect -7048 -1288 -6992 -1286
rect -6088 -1234 -6032 -1232
rect -6088 -1286 -6086 -1234
rect -6086 -1286 -6034 -1234
rect -6034 -1286 -6032 -1234
rect -6088 -1288 -6032 -1286
<< metal3 >>
rect -7200 6328 -5880 6360
rect -7200 6272 -7048 6328
rect -6992 6272 -6568 6328
rect -6512 6272 -6088 6328
rect -6032 6272 -5880 6328
rect -7200 6088 -5880 6272
rect -7200 6032 -7048 6088
rect -6992 6032 -6568 6088
rect -6512 6032 -6088 6088
rect -6032 6032 -5880 6088
rect -7200 5968 -5880 6032
rect -7200 5912 -7048 5968
rect -6992 5912 -6568 5968
rect -6512 5912 -6088 5968
rect -6032 5912 -5880 5968
rect -7200 5848 -5880 5912
rect -7200 5792 -7048 5848
rect -6992 5792 -6568 5848
rect -6512 5792 -6088 5848
rect -6032 5792 -5880 5848
rect -7200 5760 -5880 5792
rect -6600 5608 -6480 5640
rect -6600 5552 -6568 5608
rect -6512 5552 -6480 5608
rect -6600 5520 -6480 5552
rect -7200 5368 -5880 5400
rect -7200 5312 -6808 5368
rect -6752 5312 -6328 5368
rect -6272 5312 -5880 5368
rect -7200 5220 -5880 5312
rect -7200 5128 -5880 5160
rect -7200 5072 -6568 5128
rect -6512 5072 -5880 5128
rect -7200 5040 -5880 5072
rect -7200 4888 -5880 4980
rect -7200 4832 -7048 4888
rect -6992 4832 -6808 4888
rect -6752 4832 -6568 4888
rect -6512 4832 -6328 4888
rect -6272 4832 -6088 4888
rect -6032 4832 -5880 4888
rect -7200 4800 -5880 4832
rect -6840 4048 -6720 4080
rect -6840 3992 -6808 4048
rect -6752 3992 -6720 4048
rect -6840 3960 -6720 3992
rect -6360 4048 -6240 4080
rect -6360 3992 -6328 4048
rect -6272 3992 -6240 4048
rect -6360 3960 -6240 3992
rect -7200 3808 -5880 3840
rect -7200 3752 -7048 3808
rect -6992 3752 -6088 3808
rect -6032 3752 -5880 3808
rect -7200 3720 -5880 3752
rect -7200 3568 -5880 3600
rect -7200 3512 -7048 3568
rect -6992 3512 -6088 3568
rect -6032 3512 -5880 3568
rect -7200 3480 -5880 3512
rect -7200 2760 -5880 3360
rect -7200 2608 -5880 2640
rect -7200 2552 -7048 2608
rect -6992 2552 -6088 2608
rect -6032 2552 -5880 2608
rect -7200 2520 -5880 2552
rect -7200 2280 -5880 2400
rect -7200 2128 -5880 2160
rect -7200 2072 -7048 2128
rect -6992 2072 -6088 2128
rect -6032 2072 -5880 2128
rect -7200 2040 -5880 2072
rect -7200 1800 -5880 1920
rect -7200 1648 -5880 1680
rect -7200 1592 -7048 1648
rect -6992 1592 -6088 1648
rect -6032 1592 -5880 1648
rect -7200 1560 -5880 1592
rect -7200 1320 -5880 1440
rect -7200 1168 -5880 1200
rect -7200 1112 -7048 1168
rect -6992 1112 -6088 1168
rect -6032 1112 -5880 1168
rect -7200 1080 -5880 1112
rect -7200 840 -5880 960
rect -7200 688 -5880 720
rect -7200 632 -7048 688
rect -6992 632 -6088 688
rect -6032 632 -5880 688
rect -7200 600 -5880 632
rect -7200 -120 -5880 480
rect -7200 -272 -5880 -240
rect -7200 -328 -7048 -272
rect -6992 -328 -6088 -272
rect -6032 -328 -5880 -272
rect -7200 -360 -5880 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -7200 -752 -5880 -720
rect -7200 -808 -7048 -752
rect -6992 -808 -6088 -752
rect -6032 -808 -5880 -752
rect -7200 -872 -5880 -808
rect -7200 -928 -7048 -872
rect -6992 -928 -6088 -872
rect -6032 -928 -5880 -872
rect -7200 -992 -5880 -928
rect -7200 -1048 -7048 -992
rect -6992 -1048 -6088 -992
rect -6032 -1048 -5880 -992
rect -7200 -1232 -5880 -1048
rect -7200 -1288 -7048 -1232
rect -6992 -1288 -6088 -1232
rect -6032 -1288 -5880 -1232
rect -7200 -1320 -5880 -1288
<< via3 >>
rect -6568 5552 -6512 5608
rect -6808 5312 -6752 5368
rect -6328 5312 -6272 5368
rect -6568 5072 -6512 5128
rect -7048 4832 -6992 4888
rect -6808 4832 -6752 4888
rect -6328 4832 -6272 4888
rect -6088 4832 -6032 4888
rect -6808 3992 -6752 4048
rect -6328 3992 -6272 4048
rect -6808 -568 -6752 -512
rect -6328 -568 -6272 -512
<< metal4 >>
rect -6600 5608 -6480 5640
rect -6600 5552 -6568 5608
rect -6512 5552 -6480 5608
rect -6840 5368 -6720 5400
rect -6840 5312 -6808 5368
rect -6752 5312 -6720 5368
rect -7080 4888 -6960 4920
rect -7080 4832 -7048 4888
rect -6992 4832 -6960 4888
rect -7080 4800 -6960 4832
rect -6840 4888 -6720 5312
rect -6600 5128 -6480 5552
rect -6600 5072 -6568 5128
rect -6512 5072 -6480 5128
rect -6600 5040 -6480 5072
rect -6360 5368 -6240 5400
rect -6360 5312 -6328 5368
rect -6272 5312 -6240 5368
rect -6840 4832 -6808 4888
rect -6752 4832 -6720 4888
rect -6840 4800 -6720 4832
rect -6360 4888 -6240 5312
rect -6360 4832 -6328 4888
rect -6272 4832 -6240 4888
rect -6360 4800 -6240 4832
rect -6120 4888 -6000 4920
rect -6120 4832 -6088 4888
rect -6032 4832 -6000 4888
rect -6120 4800 -6000 4832
rect -6840 4048 -6720 4080
rect -6840 3992 -6808 4048
rect -6752 3992 -6720 4048
rect -6840 3840 -6720 3992
rect -7080 3720 -6720 3840
rect -6840 -512 -6720 3720
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 4048 -6240 4080
rect -6360 3992 -6328 4048
rect -6272 3992 -6240 4048
rect -6360 3840 -6240 3992
rect -6360 3720 -6000 3840
rect -6360 -512 -6240 3720
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
<< labels >>
rlabel metal1 s -6780 -900 -6780 -900 4 d1
rlabel metal1 s -6300 -900 -6300 -900 4 d2
rlabel metal1 s -6540 6540 -6540 6540 4 gnd
rlabel metal1 s -6540 5100 -6540 5100 4 gnd
rlabel metal4 s -6840 -120 -6720 3360 4 inl
port 1 nsew
rlabel metal4 s -6360 -120 -6240 3360 4 inr
port 2 nsew
rlabel metal2 s -6600 -120 -6480 3360 4 out
port 3 nsew
rlabel metal3 s -7200 5760 -5880 6360 4 vdd
port 4 nsew
rlabel metal3 s -7200 5040 -5880 5160 4 gp
port 5 nsew
rlabel metal1 s -7200 3720 -7080 3840 4 bp
port 6 nsew
rlabel metal1 s -6000 3720 -5880 3840 4 bp
port 6 nsew
rlabel metal3 s -7200 5220 -7080 5400 4 vreg
port 7 nsew
rlabel metal3 s -6000 5220 -5880 5400 4 vreg
port 7 nsew
rlabel metal3 s -7200 2760 -5880 3360 4 op
port 8 nsew
rlabel metal3 s -7200 2280 -5880 2400 4 im
port 9 nsew
rlabel metal3 s -7200 1800 -5880 1920 4 x
port 10 nsew
rlabel metal3 s -7200 1320 -5880 1440 4 y
port 11 nsew
rlabel metal3 s -7200 840 -5880 960 4 ip
port 12 nsew
rlabel metal3 s -7200 -120 -5880 480 4 om
port 13 nsew
rlabel metal3 s -7200 -1320 -5880 -720 4 gnd
port 14 nsew
<< end >>
