magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7380 4260 -6600 5460
rect -7380 2700 -6600 4020
<< nmos >>
rect -6960 -1080 -6840 -720
<< pmos >>
rect -6960 3240 -6840 3540
<< mvpmos >>
rect -6960 4800 -6840 5160
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
<< pdiff >>
rect -7080 3443 -6960 3540
rect -7080 3397 -7043 3443
rect -6997 3397 -6960 3443
rect -7080 3323 -6960 3397
rect -7080 3277 -7043 3323
rect -6997 3277 -6960 3323
rect -7080 3240 -6960 3277
rect -6840 3443 -6720 3540
rect -6840 3397 -6803 3443
rect -6757 3397 -6720 3443
rect -6840 3323 -6720 3397
rect -6840 3277 -6803 3323
rect -6757 3277 -6720 3323
rect -6840 3240 -6720 3277
<< mvpdiff >>
rect -7080 5123 -6960 5160
rect -7080 5077 -7043 5123
rect -6997 5077 -6960 5123
rect -7080 5003 -6960 5077
rect -7080 4957 -7043 5003
rect -6997 4957 -6960 5003
rect -7080 4883 -6960 4957
rect -7080 4837 -7043 4883
rect -6997 4837 -6960 4883
rect -7080 4800 -6960 4837
rect -6840 5123 -6720 5160
rect -6840 5077 -6803 5123
rect -6757 5077 -6720 5123
rect -6840 5003 -6720 5077
rect -6840 4957 -6803 5003
rect -6757 4957 -6720 5003
rect -6840 4883 -6720 4957
rect -6840 4837 -6803 4883
rect -6757 4837 -6720 4883
rect -6840 4800 -6720 4837
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
<< pdiffc >>
rect -7043 3397 -6997 3443
rect -7043 3277 -6997 3323
rect -6803 3397 -6757 3443
rect -6803 3277 -6757 3323
<< mvpdiffc >>
rect -7043 5077 -6997 5123
rect -7043 4957 -6997 5003
rect -7043 4837 -6997 4883
rect -6803 5077 -6757 5123
rect -6803 4957 -6757 5003
rect -6803 4837 -6757 4883
<< psubdiff >>
rect -7560 5603 -6600 5640
rect -7560 5557 -7523 5603
rect -7477 5557 -7403 5603
rect -7357 5557 -7283 5603
rect -7237 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6600 5603
rect -7560 5520 -6600 5557
rect -7560 5483 -7440 5520
rect -7560 5437 -7523 5483
rect -7477 5437 -7440 5483
rect -7560 5363 -7440 5437
rect -7560 5317 -7523 5363
rect -7477 5317 -7440 5363
rect -7560 5243 -7440 5317
rect -7560 5197 -7523 5243
rect -7477 5197 -7440 5243
rect -7560 5123 -7440 5197
rect -7560 5077 -7523 5123
rect -7477 5077 -7440 5123
rect -7560 5003 -7440 5077
rect -7560 4957 -7523 5003
rect -7477 4957 -7440 5003
rect -7560 4883 -7440 4957
rect -7560 4837 -7523 4883
rect -7477 4837 -7440 4883
rect -7560 4763 -7440 4837
rect -7560 4717 -7523 4763
rect -7477 4717 -7440 4763
rect -7560 4643 -7440 4717
rect -7560 4597 -7523 4643
rect -7477 4597 -7440 4643
rect -7560 4523 -7440 4597
rect -7560 4477 -7523 4523
rect -7477 4477 -7440 4523
rect -7560 4403 -7440 4477
rect -7560 4357 -7523 4403
rect -7477 4357 -7440 4403
rect -7560 4283 -7440 4357
rect -7560 4237 -7523 4283
rect -7477 4237 -7440 4283
rect -7560 4200 -7440 4237
rect -7560 4163 -6600 4200
rect -7560 4117 -7523 4163
rect -7477 4117 -7403 4163
rect -7357 4117 -7283 4163
rect -7237 4117 -7163 4163
rect -7117 4117 -7043 4163
rect -6997 4117 -6923 4163
rect -6877 4117 -6803 4163
rect -6757 4117 -6683 4163
rect -6637 4117 -6600 4163
rect -7560 4080 -6600 4117
rect -7560 4043 -7440 4080
rect -7560 3997 -7523 4043
rect -7477 3997 -7440 4043
rect -7560 3923 -7440 3997
rect -7560 3877 -7523 3923
rect -7477 3877 -7440 3923
rect -7560 3803 -7440 3877
rect -7560 3757 -7523 3803
rect -7477 3757 -7440 3803
rect -7560 3683 -7440 3757
rect -7560 3637 -7523 3683
rect -7477 3637 -7440 3683
rect -7560 3563 -7440 3637
rect -7560 3517 -7523 3563
rect -7477 3517 -7440 3563
rect -7560 3443 -7440 3517
rect -7560 3397 -7523 3443
rect -7477 3397 -7440 3443
rect -7560 3323 -7440 3397
rect -7560 3277 -7523 3323
rect -7477 3277 -7440 3323
rect -7560 3203 -7440 3277
rect -7560 3157 -7523 3203
rect -7477 3157 -7440 3203
rect -7560 3083 -7440 3157
rect -7560 3037 -7523 3083
rect -7477 3037 -7440 3083
rect -7560 2963 -7440 3037
rect -7560 2917 -7523 2963
rect -7477 2917 -7440 2963
rect -7560 2843 -7440 2917
rect -7560 2797 -7523 2843
rect -7477 2797 -7440 2843
rect -7560 2723 -7440 2797
rect -7560 2677 -7523 2723
rect -7477 2677 -7440 2723
rect -7560 2640 -7440 2677
rect -7560 2603 -6600 2640
rect -7560 2557 -7523 2603
rect -7477 2557 -7403 2603
rect -7357 2557 -7283 2603
rect -7237 2557 -7163 2603
rect -7117 2557 -7043 2603
rect -6997 2557 -6923 2603
rect -6877 2557 -6803 2603
rect -6757 2557 -6683 2603
rect -6637 2557 -6600 2603
rect -7560 2520 -6600 2557
rect -7560 2483 -7440 2520
rect -7560 2437 -7523 2483
rect -7477 2437 -7440 2483
rect -7560 2363 -7440 2437
rect -7560 2317 -7523 2363
rect -7477 2317 -7440 2363
rect -7560 2243 -7440 2317
rect -7560 2197 -7523 2243
rect -7477 2197 -7440 2243
rect -7560 2123 -7440 2197
rect -7560 2077 -7523 2123
rect -7477 2077 -7440 2123
rect -7560 2003 -7440 2077
rect -7560 1957 -7523 2003
rect -7477 1957 -7440 2003
rect -7560 1883 -7440 1957
rect -7560 1837 -7523 1883
rect -7477 1837 -7440 1883
rect -7560 1763 -7440 1837
rect -7560 1717 -7523 1763
rect -7477 1717 -7440 1763
rect -7560 1680 -7440 1717
rect -7560 1643 -6600 1680
rect -7560 1597 -7523 1643
rect -7477 1597 -7403 1643
rect -7357 1597 -7283 1643
rect -7237 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6600 1643
rect -7560 1560 -6600 1597
rect -7560 1523 -7440 1560
rect -7560 1477 -7523 1523
rect -7477 1477 -7440 1523
rect -7560 1403 -7440 1477
rect -7560 1357 -7523 1403
rect -7477 1357 -7440 1403
rect -7560 1283 -7440 1357
rect -7560 1237 -7523 1283
rect -7477 1237 -7440 1283
rect -7560 1200 -7440 1237
rect -7560 1163 -6600 1200
rect -7560 1117 -7523 1163
rect -7477 1117 -7403 1163
rect -7357 1117 -7283 1163
rect -7237 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6600 1163
rect -7560 1080 -6600 1117
rect -7560 1043 -7440 1080
rect -7560 997 -7523 1043
rect -7477 997 -7440 1043
rect -7560 923 -7440 997
rect -7560 877 -7523 923
rect -7477 877 -7440 923
rect -7560 803 -7440 877
rect -7560 757 -7523 803
rect -7477 757 -7440 803
rect -7560 720 -7440 757
rect -7560 683 -6600 720
rect -7560 637 -7523 683
rect -7477 637 -7403 683
rect -7357 637 -7283 683
rect -7237 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6600 683
rect -7560 600 -6600 637
rect -7560 563 -7440 600
rect -7560 517 -7523 563
rect -7477 517 -7440 563
rect -7560 443 -7440 517
rect -7560 397 -7523 443
rect -7477 397 -7440 443
rect -7560 323 -7440 397
rect -7560 277 -7523 323
rect -7477 277 -7440 323
rect -7560 203 -7440 277
rect -7560 157 -7523 203
rect -7477 157 -7440 203
rect -7560 83 -7440 157
rect -7560 37 -7523 83
rect -7477 37 -7440 83
rect -7560 -37 -7440 37
rect -7560 -83 -7523 -37
rect -7477 -83 -7440 -37
rect -7560 -157 -7440 -83
rect -7560 -203 -7523 -157
rect -7477 -203 -7440 -157
rect -7560 -240 -7440 -203
rect -7560 -277 -6600 -240
rect -7560 -323 -7523 -277
rect -7477 -323 -7403 -277
rect -7357 -323 -7283 -277
rect -7237 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6600 -277
rect -7560 -360 -6600 -323
rect -7560 -397 -7440 -360
rect -7560 -443 -7523 -397
rect -7477 -443 -7440 -397
rect -7560 -517 -7440 -443
rect -7560 -563 -7523 -517
rect -7477 -563 -7440 -517
rect -7560 -637 -7440 -563
rect -7560 -683 -7523 -637
rect -7477 -683 -7440 -637
rect -7560 -757 -7440 -683
rect -7560 -803 -7523 -757
rect -7477 -803 -7440 -757
rect -7560 -877 -7440 -803
rect -7560 -923 -7523 -877
rect -7477 -923 -7440 -877
rect -7560 -997 -7440 -923
rect -7560 -1043 -7523 -997
rect -7477 -1043 -7440 -997
rect -7560 -1117 -7440 -1043
rect -7560 -1163 -7523 -1117
rect -7477 -1163 -7440 -1117
rect -7560 -1200 -7440 -1163
rect -7560 -1237 -6600 -1200
rect -7560 -1283 -7523 -1237
rect -7477 -1283 -7403 -1237
rect -7357 -1283 -7283 -1237
rect -7237 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6600 -1237
rect -7560 -1320 -6600 -1283
<< nsubdiff >>
rect -7320 3923 -6720 3960
rect -7320 3877 -7283 3923
rect -7237 3877 -7163 3923
rect -7117 3877 -7043 3923
rect -6997 3877 -6923 3923
rect -6877 3877 -6803 3923
rect -6757 3877 -6720 3923
rect -7320 3840 -6720 3877
rect -7320 3803 -7200 3840
rect -7320 3757 -7283 3803
rect -7237 3757 -7200 3803
rect -7320 3683 -7200 3757
rect -7320 3637 -7283 3683
rect -7237 3637 -7200 3683
rect -7320 3563 -7200 3637
rect -7320 3517 -7283 3563
rect -7237 3517 -7200 3563
rect -7320 3443 -7200 3517
rect -7320 3397 -7283 3443
rect -7237 3397 -7200 3443
rect -7320 3323 -7200 3397
rect -7320 3277 -7283 3323
rect -7237 3277 -7200 3323
rect -7320 3203 -7200 3277
rect -7320 3157 -7283 3203
rect -7237 3157 -7200 3203
rect -7320 3083 -7200 3157
rect -7320 3037 -7283 3083
rect -7237 3037 -7200 3083
rect -7320 2963 -7200 3037
rect -7320 2917 -7283 2963
rect -7237 2917 -7200 2963
rect -7320 2880 -7200 2917
rect -7320 2843 -6720 2880
rect -7320 2797 -7283 2843
rect -7237 2797 -7163 2843
rect -7117 2797 -7043 2843
rect -6997 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6720 2843
rect -7320 2760 -6720 2797
<< mvnsubdiff >>
rect -7320 5363 -6720 5400
rect -7320 5317 -7283 5363
rect -7237 5317 -7163 5363
rect -7117 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6720 5363
rect -7320 5280 -6720 5317
rect -7320 5243 -7200 5280
rect -7320 5197 -7283 5243
rect -7237 5197 -7200 5243
rect -7320 5123 -7200 5197
rect -7320 5077 -7283 5123
rect -7237 5077 -7200 5123
rect -7320 5003 -7200 5077
rect -7320 4957 -7283 5003
rect -7237 4957 -7200 5003
rect -7320 4883 -7200 4957
rect -7320 4837 -7283 4883
rect -7237 4837 -7200 4883
rect -7320 4763 -7200 4837
rect -7320 4717 -7283 4763
rect -7237 4717 -7200 4763
rect -7320 4643 -7200 4717
rect -7320 4597 -7283 4643
rect -7237 4597 -7200 4643
rect -7320 4523 -7200 4597
rect -7320 4477 -7283 4523
rect -7237 4477 -7200 4523
rect -7320 4440 -7200 4477
rect -7320 4403 -6720 4440
rect -7320 4357 -7283 4403
rect -7237 4357 -7163 4403
rect -7117 4357 -7043 4403
rect -6997 4357 -6923 4403
rect -6877 4357 -6803 4403
rect -6757 4357 -6720 4403
rect -7320 4320 -6720 4357
<< psubdiffcont >>
rect -7523 5557 -7477 5603
rect -7403 5557 -7357 5603
rect -7283 5557 -7237 5603
rect -7163 5557 -7117 5603
rect -7043 5557 -6997 5603
rect -6923 5557 -6877 5603
rect -6803 5557 -6757 5603
rect -6683 5557 -6637 5603
rect -7523 5437 -7477 5483
rect -7523 5317 -7477 5363
rect -7523 5197 -7477 5243
rect -7523 5077 -7477 5123
rect -7523 4957 -7477 5003
rect -7523 4837 -7477 4883
rect -7523 4717 -7477 4763
rect -7523 4597 -7477 4643
rect -7523 4477 -7477 4523
rect -7523 4357 -7477 4403
rect -7523 4237 -7477 4283
rect -7523 4117 -7477 4163
rect -7403 4117 -7357 4163
rect -7283 4117 -7237 4163
rect -7163 4117 -7117 4163
rect -7043 4117 -6997 4163
rect -6923 4117 -6877 4163
rect -6803 4117 -6757 4163
rect -6683 4117 -6637 4163
rect -7523 3997 -7477 4043
rect -7523 3877 -7477 3923
rect -7523 3757 -7477 3803
rect -7523 3637 -7477 3683
rect -7523 3517 -7477 3563
rect -7523 3397 -7477 3443
rect -7523 3277 -7477 3323
rect -7523 3157 -7477 3203
rect -7523 3037 -7477 3083
rect -7523 2917 -7477 2963
rect -7523 2797 -7477 2843
rect -7523 2677 -7477 2723
rect -7523 2557 -7477 2603
rect -7403 2557 -7357 2603
rect -7283 2557 -7237 2603
rect -7163 2557 -7117 2603
rect -7043 2557 -6997 2603
rect -6923 2557 -6877 2603
rect -6803 2557 -6757 2603
rect -6683 2557 -6637 2603
rect -7523 2437 -7477 2483
rect -7523 2317 -7477 2363
rect -7523 2197 -7477 2243
rect -7523 2077 -7477 2123
rect -7523 1957 -7477 2003
rect -7523 1837 -7477 1883
rect -7523 1717 -7477 1763
rect -7523 1597 -7477 1643
rect -7403 1597 -7357 1643
rect -7283 1597 -7237 1643
rect -7163 1597 -7117 1643
rect -7043 1597 -6997 1643
rect -6923 1597 -6877 1643
rect -6803 1597 -6757 1643
rect -6683 1597 -6637 1643
rect -7523 1477 -7477 1523
rect -7523 1357 -7477 1403
rect -7523 1237 -7477 1283
rect -7523 1117 -7477 1163
rect -7403 1117 -7357 1163
rect -7283 1117 -7237 1163
rect -7163 1117 -7117 1163
rect -7043 1117 -6997 1163
rect -6923 1117 -6877 1163
rect -6803 1117 -6757 1163
rect -6683 1117 -6637 1163
rect -7523 997 -7477 1043
rect -7523 877 -7477 923
rect -7523 757 -7477 803
rect -7523 637 -7477 683
rect -7403 637 -7357 683
rect -7283 637 -7237 683
rect -7163 637 -7117 683
rect -7043 637 -6997 683
rect -6923 637 -6877 683
rect -6803 637 -6757 683
rect -6683 637 -6637 683
rect -7523 517 -7477 563
rect -7523 397 -7477 443
rect -7523 277 -7477 323
rect -7523 157 -7477 203
rect -7523 37 -7477 83
rect -7523 -83 -7477 -37
rect -7523 -203 -7477 -157
rect -7523 -323 -7477 -277
rect -7403 -323 -7357 -277
rect -7283 -323 -7237 -277
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -7523 -443 -7477 -397
rect -7523 -563 -7477 -517
rect -7523 -683 -7477 -637
rect -7523 -803 -7477 -757
rect -7523 -923 -7477 -877
rect -7523 -1043 -7477 -997
rect -7523 -1163 -7477 -1117
rect -7523 -1283 -7477 -1237
rect -7403 -1283 -7357 -1237
rect -7283 -1283 -7237 -1237
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
<< nsubdiffcont >>
rect -7283 3877 -7237 3923
rect -7163 3877 -7117 3923
rect -7043 3877 -6997 3923
rect -6923 3877 -6877 3923
rect -6803 3877 -6757 3923
rect -7283 3757 -7237 3803
rect -7283 3637 -7237 3683
rect -7283 3517 -7237 3563
rect -7283 3397 -7237 3443
rect -7283 3277 -7237 3323
rect -7283 3157 -7237 3203
rect -7283 3037 -7237 3083
rect -7283 2917 -7237 2963
rect -7283 2797 -7237 2843
rect -7163 2797 -7117 2843
rect -7043 2797 -6997 2843
rect -6923 2797 -6877 2843
rect -6803 2797 -6757 2843
<< mvnsubdiffcont >>
rect -7283 5317 -7237 5363
rect -7163 5317 -7117 5363
rect -7043 5317 -6997 5363
rect -6923 5317 -6877 5363
rect -6803 5317 -6757 5363
rect -7283 5197 -7237 5243
rect -7283 5077 -7237 5123
rect -7283 4957 -7237 5003
rect -7283 4837 -7237 4883
rect -7283 4717 -7237 4763
rect -7283 4597 -7237 4643
rect -7283 4477 -7237 4523
rect -7283 4357 -7237 4403
rect -7163 4357 -7117 4403
rect -7043 4357 -6997 4403
rect -6923 4357 -6877 4403
rect -6803 4357 -6757 4403
<< polysilicon >>
rect -6960 5160 -6840 5220
rect -6960 4643 -6840 4800
rect -6960 4597 -6923 4643
rect -6877 4597 -6840 4643
rect -6960 4560 -6840 4597
rect -6960 3540 -6840 3600
rect -6960 3083 -6840 3240
rect -6960 3037 -6923 3083
rect -6877 3037 -6840 3083
rect -6960 3000 -6840 3037
rect -6960 -517 -6840 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6840 -517
rect -6960 -720 -6840 -563
rect -6960 -1140 -6840 -1080
<< polycontact >>
rect -6923 4597 -6877 4643
rect -6923 3037 -6877 3083
rect -6923 -563 -6877 -517
<< metal1 >>
rect -7560 5603 -6600 5640
rect -7560 5557 -7523 5603
rect -7477 5557 -7403 5603
rect -7357 5557 -7283 5603
rect -7237 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6600 5603
rect -7560 5520 -6600 5557
rect -7560 5483 -7440 5520
rect -7560 5437 -7523 5483
rect -7477 5437 -7440 5483
rect -7560 5363 -7440 5437
rect -7560 5317 -7523 5363
rect -7477 5317 -7440 5363
rect -7560 5243 -7440 5317
rect -7560 5197 -7523 5243
rect -7477 5197 -7440 5243
rect -7560 5123 -7440 5197
rect -7560 5077 -7523 5123
rect -7477 5077 -7440 5123
rect -7560 5003 -7440 5077
rect -7560 4957 -7523 5003
rect -7477 4957 -7440 5003
rect -7560 4883 -7440 4957
rect -7560 4837 -7523 4883
rect -7477 4837 -7440 4883
rect -7560 4763 -7440 4837
rect -7560 4717 -7523 4763
rect -7477 4717 -7440 4763
rect -7560 4643 -7440 4717
rect -7560 4597 -7523 4643
rect -7477 4597 -7440 4643
rect -7560 4523 -7440 4597
rect -7560 4477 -7523 4523
rect -7477 4477 -7440 4523
rect -7560 4403 -7440 4477
rect -7560 4357 -7523 4403
rect -7477 4357 -7440 4403
rect -7560 4283 -7440 4357
rect -7320 5366 -6600 5400
rect -7320 5363 -6806 5366
rect -7320 5317 -7283 5363
rect -7237 5317 -7163 5363
rect -7117 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6806 5363
rect -7320 5314 -6806 5317
rect -6754 5314 -6600 5366
rect -7320 5280 -6600 5314
rect -7320 5243 -7200 5280
rect -7320 5197 -7283 5243
rect -7237 5197 -7200 5243
rect -7320 5123 -7200 5197
rect -7320 5077 -7283 5123
rect -7237 5077 -7200 5123
rect -7320 5003 -7200 5077
rect -7320 4957 -7283 5003
rect -7237 4957 -7200 5003
rect -7320 4883 -7200 4957
rect -7320 4837 -7283 4883
rect -7237 4837 -7200 4883
rect -7320 4763 -7200 4837
rect -7320 4717 -7283 4763
rect -7237 4717 -7200 4763
rect -7320 4643 -7200 4717
rect -7320 4597 -7283 4643
rect -7237 4597 -7200 4643
rect -7320 4523 -7200 4597
rect -7080 5123 -6960 5160
rect -7080 5077 -7043 5123
rect -6997 5077 -6960 5123
rect -7080 5003 -6960 5077
rect -7080 4957 -7043 5003
rect -6997 4957 -6960 5003
rect -7080 4883 -6960 4957
rect -7080 4837 -7043 4883
rect -6997 4837 -6960 4883
rect -7080 4680 -6960 4837
rect -6840 5126 -6720 5160
rect -6840 5074 -6806 5126
rect -6754 5074 -6720 5126
rect -6840 5006 -6720 5074
rect -6840 4954 -6806 5006
rect -6754 4954 -6720 5006
rect -6840 4886 -6720 4954
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4800 -6720 4834
rect -7080 4643 -6840 4680
rect -7080 4597 -6923 4643
rect -6877 4597 -6840 4643
rect -7080 4560 -6840 4597
rect -7320 4477 -7283 4523
rect -7237 4477 -7200 4523
rect -7320 4440 -7200 4477
rect -7320 4403 -6600 4440
rect -7320 4357 -7283 4403
rect -7237 4357 -7163 4403
rect -7117 4357 -7043 4403
rect -6997 4357 -6923 4403
rect -6877 4357 -6803 4403
rect -6757 4357 -6600 4403
rect -7320 4320 -6600 4357
rect -7560 4237 -7523 4283
rect -7477 4237 -7440 4283
rect -7560 4200 -7440 4237
rect -7560 4163 -6600 4200
rect -7560 4117 -7523 4163
rect -7477 4117 -7403 4163
rect -7357 4117 -7283 4163
rect -7237 4117 -7163 4163
rect -7117 4117 -7043 4163
rect -6997 4117 -6923 4163
rect -6877 4117 -6803 4163
rect -6757 4117 -6683 4163
rect -6637 4117 -6600 4163
rect -7560 4080 -6600 4117
rect -7560 4043 -7440 4080
rect -7560 3997 -7523 4043
rect -7477 3997 -7440 4043
rect -7560 3923 -7440 3997
rect -7560 3877 -7523 3923
rect -7477 3877 -7440 3923
rect -7560 3803 -7440 3877
rect -7560 3757 -7523 3803
rect -7477 3757 -7440 3803
rect -7560 3683 -7440 3757
rect -7560 3637 -7523 3683
rect -7477 3637 -7440 3683
rect -7560 3563 -7440 3637
rect -7560 3517 -7523 3563
rect -7477 3517 -7440 3563
rect -7560 3443 -7440 3517
rect -7560 3397 -7523 3443
rect -7477 3397 -7440 3443
rect -7560 3323 -7440 3397
rect -7560 3277 -7523 3323
rect -7477 3277 -7440 3323
rect -7560 3203 -7440 3277
rect -7560 3157 -7523 3203
rect -7477 3157 -7440 3203
rect -7560 3083 -7440 3157
rect -7560 3037 -7523 3083
rect -7477 3037 -7440 3083
rect -7560 2963 -7440 3037
rect -7560 2917 -7523 2963
rect -7477 2917 -7440 2963
rect -7560 2843 -7440 2917
rect -7560 2797 -7523 2843
rect -7477 2797 -7440 2843
rect -7560 2723 -7440 2797
rect -7320 3923 -6720 3960
rect -7320 3877 -7283 3923
rect -7237 3877 -7163 3923
rect -7117 3877 -7043 3923
rect -6997 3877 -6923 3923
rect -6877 3877 -6803 3923
rect -6757 3877 -6720 3923
rect -7320 3840 -6720 3877
rect -7320 3803 -7200 3840
rect -7320 3757 -7283 3803
rect -7237 3757 -7200 3803
rect -7320 3683 -7200 3757
rect -7320 3637 -7283 3683
rect -7237 3637 -7200 3683
rect -7320 3563 -7200 3637
rect -7320 3517 -7283 3563
rect -7237 3517 -7200 3563
rect -7320 3443 -7200 3517
rect -7320 3397 -7283 3443
rect -7237 3397 -7200 3443
rect -7320 3323 -7200 3397
rect -7320 3277 -7283 3323
rect -7237 3277 -7200 3323
rect -7320 3203 -7200 3277
rect -7320 3157 -7283 3203
rect -7237 3157 -7200 3203
rect -7320 3083 -7200 3157
rect -7320 3037 -7283 3083
rect -7237 3037 -7200 3083
rect -7320 2963 -7200 3037
rect -7080 3443 -6960 3540
rect -7080 3397 -7043 3443
rect -6997 3397 -6960 3443
rect -7080 3323 -6960 3397
rect -7080 3277 -7043 3323
rect -6997 3277 -6960 3323
rect -7080 3120 -6960 3277
rect -6840 3446 -6720 3540
rect -6840 3394 -6806 3446
rect -6754 3394 -6720 3446
rect -6840 3326 -6720 3394
rect -6840 3274 -6806 3326
rect -6754 3274 -6720 3326
rect -6840 3240 -6720 3274
rect -7080 3083 -6840 3120
rect -7080 3037 -6923 3083
rect -6877 3037 -6840 3083
rect -7080 3000 -6840 3037
rect -7320 2917 -7283 2963
rect -7237 2917 -7200 2963
rect -7320 2880 -7200 2917
rect -7320 2846 -6600 2880
rect -7320 2794 -7286 2846
rect -7234 2843 -6600 2846
rect -7234 2797 -7163 2843
rect -7117 2797 -7043 2843
rect -6997 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6600 2843
rect -7234 2794 -6600 2797
rect -7320 2760 -6600 2794
rect -7560 2677 -7523 2723
rect -7477 2677 -7440 2723
rect -7560 2640 -7440 2677
rect -7560 2606 -6600 2640
rect -7560 2603 -6806 2606
rect -6754 2603 -6600 2606
rect -7560 2557 -7523 2603
rect -7477 2557 -7403 2603
rect -7357 2557 -7283 2603
rect -7237 2557 -7163 2603
rect -7117 2557 -7043 2603
rect -6997 2557 -6923 2603
rect -6877 2557 -6806 2603
rect -6754 2557 -6683 2603
rect -6637 2557 -6600 2603
rect -7560 2554 -6806 2557
rect -6754 2554 -6600 2557
rect -7560 2520 -6600 2554
rect -7560 2483 -7440 2520
rect -7560 2437 -7523 2483
rect -7477 2437 -7440 2483
rect -7560 2363 -7440 2437
rect -7560 2317 -7523 2363
rect -7477 2317 -7440 2363
rect -7560 2243 -7440 2317
rect -7560 2197 -7523 2243
rect -7477 2197 -7440 2243
rect -7560 2123 -7440 2197
rect -7560 2077 -7523 2123
rect -7477 2077 -7440 2123
rect -7560 2003 -7440 2077
rect -7560 1957 -7523 2003
rect -7477 1957 -7440 2003
rect -7560 1883 -7440 1957
rect -7560 1837 -7523 1883
rect -7477 1837 -7440 1883
rect -7560 1763 -7440 1837
rect -7560 1717 -7523 1763
rect -7477 1717 -7440 1763
rect -7560 1680 -7440 1717
rect -7560 1646 -6600 1680
rect -7560 1643 -6806 1646
rect -6754 1643 -6600 1646
rect -7560 1597 -7523 1643
rect -7477 1597 -7403 1643
rect -7357 1597 -7283 1643
rect -7237 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6806 1643
rect -6754 1597 -6683 1643
rect -6637 1597 -6600 1643
rect -7560 1594 -6806 1597
rect -6754 1594 -6600 1597
rect -7560 1560 -6600 1594
rect -7560 1523 -7440 1560
rect -7560 1477 -7523 1523
rect -7477 1477 -7440 1523
rect -7560 1403 -7440 1477
rect -7560 1357 -7523 1403
rect -7477 1357 -7440 1403
rect -7560 1283 -7440 1357
rect -7560 1237 -7523 1283
rect -7477 1237 -7440 1283
rect -7560 1200 -7440 1237
rect -7560 1166 -6600 1200
rect -7560 1163 -6806 1166
rect -6754 1163 -6600 1166
rect -7560 1117 -7523 1163
rect -7477 1117 -7403 1163
rect -7357 1117 -7283 1163
rect -7237 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6806 1163
rect -6754 1117 -6683 1163
rect -6637 1117 -6600 1163
rect -7560 1114 -6806 1117
rect -6754 1114 -6600 1117
rect -7560 1080 -6600 1114
rect -7560 1043 -7440 1080
rect -7560 997 -7523 1043
rect -7477 997 -7440 1043
rect -7560 923 -7440 997
rect -7560 877 -7523 923
rect -7477 877 -7440 923
rect -7560 803 -7440 877
rect -7560 757 -7523 803
rect -7477 757 -7440 803
rect -7560 720 -7440 757
rect -7560 686 -6600 720
rect -7560 683 -6806 686
rect -6754 683 -6600 686
rect -7560 637 -7523 683
rect -7477 637 -7403 683
rect -7357 637 -7283 683
rect -7237 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6806 683
rect -6754 637 -6683 683
rect -6637 637 -6600 683
rect -7560 634 -6806 637
rect -6754 634 -6600 637
rect -7560 600 -6600 634
rect -7560 563 -7440 600
rect -7560 517 -7523 563
rect -7477 517 -7440 563
rect -7560 443 -7440 517
rect -7560 397 -7523 443
rect -7477 397 -7440 443
rect -7560 323 -7440 397
rect -7560 277 -7523 323
rect -7477 277 -7440 323
rect -7560 203 -7440 277
rect -7560 157 -7523 203
rect -7477 157 -7440 203
rect -7560 83 -7440 157
rect -7560 37 -7523 83
rect -7477 37 -7440 83
rect -7560 -37 -7440 37
rect -7560 -83 -7523 -37
rect -7477 -83 -7440 -37
rect -7560 -157 -7440 -83
rect -7560 -203 -7523 -157
rect -7477 -203 -7440 -157
rect -7560 -240 -7440 -203
rect -7560 -274 -6600 -240
rect -7560 -277 -6806 -274
rect -6754 -277 -6600 -274
rect -7560 -323 -7523 -277
rect -7477 -323 -7403 -277
rect -7357 -323 -7283 -277
rect -7237 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6806 -277
rect -6754 -323 -6683 -277
rect -6637 -323 -6600 -277
rect -7560 -326 -6806 -323
rect -6754 -326 -6600 -323
rect -7560 -360 -6600 -326
rect -7560 -397 -7440 -360
rect -7560 -443 -7523 -397
rect -7477 -443 -7440 -397
rect -7560 -517 -7440 -443
rect -7560 -563 -7523 -517
rect -7477 -563 -7440 -517
rect -7560 -637 -7440 -563
rect -7560 -683 -7523 -637
rect -7477 -683 -7440 -637
rect -7560 -757 -7440 -683
rect -7560 -803 -7523 -757
rect -7477 -803 -7440 -757
rect -7560 -877 -7440 -803
rect -7560 -923 -7523 -877
rect -7477 -923 -7440 -877
rect -7560 -997 -7440 -923
rect -7560 -1043 -7523 -997
rect -7477 -1043 -7440 -997
rect -7560 -1117 -7440 -1043
rect -7080 -517 -6840 -480
rect -7080 -563 -6923 -517
rect -6877 -563 -6840 -517
rect -7080 -600 -6840 -563
rect -7080 -757 -6960 -600
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -754 -6720 -720
rect -6840 -806 -6806 -754
rect -6754 -806 -6720 -754
rect -6840 -874 -6720 -806
rect -6840 -926 -6806 -874
rect -6754 -926 -6720 -874
rect -6840 -994 -6720 -926
rect -6840 -1046 -6806 -994
rect -6754 -1046 -6720 -994
rect -6840 -1080 -6720 -1046
rect -7560 -1163 -7523 -1117
rect -7477 -1163 -7440 -1117
rect -7560 -1200 -7440 -1163
rect -7560 -1234 -6600 -1200
rect -7560 -1237 -6806 -1234
rect -6754 -1237 -6600 -1234
rect -7560 -1283 -7523 -1237
rect -7477 -1283 -7403 -1237
rect -7357 -1283 -7283 -1237
rect -7237 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6806 -1237
rect -6754 -1283 -6683 -1237
rect -6637 -1283 -6600 -1237
rect -7560 -1286 -6806 -1283
rect -6754 -1286 -6600 -1283
rect -7560 -1320 -6600 -1286
<< via1 >>
rect -6806 5363 -6754 5366
rect -6806 5317 -6803 5363
rect -6803 5317 -6757 5363
rect -6757 5317 -6754 5363
rect -6806 5314 -6754 5317
rect -6806 5123 -6754 5126
rect -6806 5077 -6803 5123
rect -6803 5077 -6757 5123
rect -6757 5077 -6754 5123
rect -6806 5074 -6754 5077
rect -6806 5003 -6754 5006
rect -6806 4957 -6803 5003
rect -6803 4957 -6757 5003
rect -6757 4957 -6754 5003
rect -6806 4954 -6754 4957
rect -6806 4883 -6754 4886
rect -6806 4837 -6803 4883
rect -6803 4837 -6757 4883
rect -6757 4837 -6754 4883
rect -6806 4834 -6754 4837
rect -6806 3443 -6754 3446
rect -6806 3397 -6803 3443
rect -6803 3397 -6757 3443
rect -6757 3397 -6754 3443
rect -6806 3394 -6754 3397
rect -6806 3323 -6754 3326
rect -6806 3277 -6803 3323
rect -6803 3277 -6757 3323
rect -6757 3277 -6754 3323
rect -6806 3274 -6754 3277
rect -7286 2843 -7234 2846
rect -7286 2797 -7283 2843
rect -7283 2797 -7237 2843
rect -7237 2797 -7234 2843
rect -7286 2794 -7234 2797
rect -6806 2603 -6754 2606
rect -6806 2557 -6803 2603
rect -6803 2557 -6757 2603
rect -6757 2557 -6754 2603
rect -6806 2554 -6754 2557
rect -6806 1643 -6754 1646
rect -6806 1597 -6803 1643
rect -6803 1597 -6757 1643
rect -6757 1597 -6754 1643
rect -6806 1594 -6754 1597
rect -6806 1163 -6754 1166
rect -6806 1117 -6803 1163
rect -6803 1117 -6757 1163
rect -6757 1117 -6754 1163
rect -6806 1114 -6754 1117
rect -6806 683 -6754 686
rect -6806 637 -6803 683
rect -6803 637 -6757 683
rect -6757 637 -6754 683
rect -6806 634 -6754 637
rect -6806 -277 -6754 -274
rect -6806 -323 -6803 -277
rect -6803 -323 -6757 -277
rect -6757 -323 -6754 -277
rect -6806 -326 -6754 -323
rect -6806 -757 -6754 -754
rect -6806 -803 -6803 -757
rect -6803 -803 -6757 -757
rect -6757 -803 -6754 -757
rect -6806 -806 -6754 -803
rect -6806 -877 -6754 -874
rect -6806 -923 -6803 -877
rect -6803 -923 -6757 -877
rect -6757 -923 -6754 -877
rect -6806 -926 -6754 -923
rect -6806 -997 -6754 -994
rect -6806 -1043 -6803 -997
rect -6803 -1043 -6757 -997
rect -6757 -1043 -6754 -997
rect -6806 -1046 -6754 -1043
rect -6806 -1237 -6754 -1234
rect -6806 -1283 -6803 -1237
rect -6803 -1283 -6757 -1237
rect -6757 -1283 -6754 -1237
rect -6806 -1286 -6754 -1283
<< metal2 >>
rect -6840 5368 -6720 5400
rect -6840 5312 -6808 5368
rect -6752 5312 -6720 5368
rect -6840 5128 -6720 5312
rect -6840 5072 -6808 5128
rect -6752 5072 -6720 5128
rect -6840 5008 -6720 5072
rect -6840 4952 -6808 5008
rect -6752 4952 -6720 5008
rect -6840 4888 -6720 4952
rect -6840 4832 -6808 4888
rect -6752 4832 -6720 4888
rect -6840 4800 -6720 4832
rect -7080 4408 -6960 4440
rect -7080 4352 -7048 4408
rect -6992 4352 -6960 4408
rect -7080 3928 -6960 4352
rect -7080 3872 -7048 3928
rect -6992 3872 -6960 3928
rect -7080 3840 -6960 3872
rect -6840 3928 -6720 3960
rect -6840 3872 -6808 3928
rect -6752 3872 -6720 3928
rect -6840 3446 -6720 3872
rect -6840 3394 -6806 3446
rect -6754 3394 -6720 3446
rect -6840 3326 -6720 3394
rect -6840 3274 -6806 3326
rect -6754 3274 -6720 3326
rect -6840 3240 -6720 3274
rect -7320 2848 -7200 2880
rect -7320 2792 -7288 2848
rect -7232 2792 -7200 2848
rect -7320 2760 -7200 2792
rect -6840 2608 -6720 2640
rect -6840 2552 -6808 2608
rect -6752 2552 -6720 2608
rect -6840 1648 -6720 2552
rect -6840 1592 -6808 1648
rect -6752 1592 -6720 1648
rect -6840 1168 -6720 1592
rect -6840 1112 -6808 1168
rect -6752 1112 -6720 1168
rect -6840 688 -6720 1112
rect -6840 632 -6808 688
rect -6752 632 -6720 688
rect -6840 -272 -6720 632
rect -6840 -328 -6808 -272
rect -6752 -328 -6720 -272
rect -6840 -754 -6720 -328
rect -6840 -806 -6806 -754
rect -6754 -806 -6720 -754
rect -6840 -874 -6720 -806
rect -6840 -926 -6806 -874
rect -6754 -926 -6720 -874
rect -6840 -994 -6720 -926
rect -6840 -1046 -6806 -994
rect -6754 -1046 -6720 -994
rect -6840 -1232 -6720 -1046
rect -6840 -1288 -6808 -1232
rect -6752 -1288 -6720 -1232
rect -6840 -1320 -6720 -1288
<< via2 >>
rect -6808 5366 -6752 5368
rect -6808 5314 -6806 5366
rect -6806 5314 -6754 5366
rect -6754 5314 -6752 5366
rect -6808 5312 -6752 5314
rect -6808 5126 -6752 5128
rect -6808 5074 -6806 5126
rect -6806 5074 -6754 5126
rect -6754 5074 -6752 5126
rect -6808 5072 -6752 5074
rect -6808 5006 -6752 5008
rect -6808 4954 -6806 5006
rect -6806 4954 -6754 5006
rect -6754 4954 -6752 5006
rect -6808 4952 -6752 4954
rect -6808 4886 -6752 4888
rect -6808 4834 -6806 4886
rect -6806 4834 -6754 4886
rect -6754 4834 -6752 4886
rect -6808 4832 -6752 4834
rect -7048 4352 -6992 4408
rect -7048 3872 -6992 3928
rect -6808 3872 -6752 3928
rect -7288 2846 -7232 2848
rect -7288 2794 -7286 2846
rect -7286 2794 -7234 2846
rect -7234 2794 -7232 2846
rect -7288 2792 -7232 2794
rect -6808 2606 -6752 2608
rect -6808 2554 -6806 2606
rect -6806 2554 -6754 2606
rect -6754 2554 -6752 2606
rect -6808 2552 -6752 2554
rect -6808 1646 -6752 1648
rect -6808 1594 -6806 1646
rect -6806 1594 -6754 1646
rect -6754 1594 -6752 1646
rect -6808 1592 -6752 1594
rect -6808 1166 -6752 1168
rect -6808 1114 -6806 1166
rect -6806 1114 -6754 1166
rect -6754 1114 -6752 1166
rect -6808 1112 -6752 1114
rect -6808 686 -6752 688
rect -6808 634 -6806 686
rect -6806 634 -6754 686
rect -6754 634 -6752 686
rect -6808 632 -6752 634
rect -6808 -274 -6752 -272
rect -6808 -326 -6806 -274
rect -6806 -326 -6754 -274
rect -6754 -326 -6752 -274
rect -6808 -328 -6752 -326
rect -6808 -1234 -6752 -1232
rect -6808 -1286 -6806 -1234
rect -6806 -1286 -6754 -1234
rect -6754 -1286 -6752 -1234
rect -6808 -1288 -6752 -1286
<< metal3 >>
rect -7560 5368 -6600 5400
rect -7560 5312 -6808 5368
rect -6752 5312 -6600 5368
rect -7560 5128 -6600 5312
rect -7560 5072 -6808 5128
rect -6752 5072 -6600 5128
rect -7560 5008 -6600 5072
rect -7560 4952 -6808 5008
rect -6752 4952 -6600 5008
rect -7560 4888 -6600 4952
rect -7560 4832 -6808 4888
rect -6752 4832 -6600 4888
rect -7560 4800 -6600 4832
rect -7560 4408 -6600 4440
rect -7560 4352 -7048 4408
rect -6992 4352 -6600 4408
rect -7560 4260 -6600 4352
rect -7560 4080 -6600 4200
rect -7560 3928 -6600 4020
rect -7560 3872 -7048 3928
rect -6992 3872 -6808 3928
rect -6752 3872 -6600 3928
rect -7560 3840 -6600 3872
rect -7560 2848 -6600 2880
rect -7560 2792 -7288 2848
rect -7232 2792 -6600 2848
rect -7560 2760 -6600 2792
rect -7560 2608 -6600 2640
rect -7560 2552 -6808 2608
rect -6752 2552 -6600 2608
rect -7560 2520 -6600 2552
rect -7560 1800 -6600 2400
rect -7560 1648 -6600 1680
rect -7560 1592 -6808 1648
rect -6752 1592 -6600 1648
rect -7560 1560 -6600 1592
rect -7560 1320 -6600 1440
rect -7560 1168 -6600 1200
rect -7560 1112 -6808 1168
rect -6752 1112 -6600 1168
rect -7560 1080 -6600 1112
rect -7560 840 -6600 960
rect -7560 688 -6600 720
rect -7560 632 -6808 688
rect -6752 632 -6600 688
rect -7560 600 -6600 632
rect -7560 -120 -6600 480
rect -7560 -272 -6600 -240
rect -7560 -328 -6808 -272
rect -6752 -328 -6600 -272
rect -7560 -360 -6600 -328
rect -7560 -1232 -6600 -720
rect -7560 -1288 -6808 -1232
rect -6752 -1288 -6600 -1232
rect -7560 -1320 -6600 -1288
<< labels >>
rlabel metal1 s -7020 4620 -7020 4620 4 hih
rlabel metal1 s -7020 3060 -7020 3060 4 hi
rlabel metal1 s -7020 -540 -7020 -540 4 lo
rlabel metal3 s -7560 4800 -6600 5400 4 vdd
port 1 nsew
rlabel metal3 s -7560 4080 -6600 4200 4 gp
port 2 nsew
rlabel metal3 s -7560 2760 -6600 2880 4 bp
port 3 nsew
rlabel metal3 s -7560 4320 -6600 4440 4 vreg
port 4 nsew
rlabel metal3 s -7560 1800 -6600 2400 4 op
port 5 nsew
rlabel metal3 s -7560 1320 -6600 1440 4 im
port 6 nsew
rlabel metal3 s -7560 840 -6600 960 4 ip
port 7 nsew
rlabel metal3 s -7560 -120 -6600 480 4 om
port 8 nsew
rlabel metal3 s -7560 -1320 -6600 -720 4 gnd
port 9 nsew
<< end >>
