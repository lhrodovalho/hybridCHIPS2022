magic
tech gf180mcuC
timestamp 1664998004
<< nwell >>
rect -738 570 -660 690
rect -738 414 -660 546
<< nmos >>
rect -696 -108 -684 -72
<< pmos >>
rect -696 468 -684 498
<< mvpmos >>
rect -696 624 -684 660
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
<< pdiff >>
rect -708 489 -696 498
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 477 -696 483
rect -708 471 -705 477
rect -699 471 -696 477
rect -708 468 -696 471
rect -684 489 -672 498
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 477 -672 483
rect -684 471 -681 477
rect -675 471 -672 477
rect -684 468 -672 471
<< mvpdiff >>
rect -708 657 -696 660
rect -708 651 -705 657
rect -699 651 -696 657
rect -708 645 -696 651
rect -708 639 -705 645
rect -699 639 -696 645
rect -708 633 -696 639
rect -708 627 -705 633
rect -699 627 -696 633
rect -708 624 -696 627
rect -684 657 -672 660
rect -684 651 -681 657
rect -675 651 -672 657
rect -684 645 -672 651
rect -684 639 -681 645
rect -675 639 -672 645
rect -684 633 -672 639
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 624 -672 627
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
<< pdiffc >>
rect -705 483 -699 489
rect -705 471 -699 477
rect -681 483 -675 489
rect -681 471 -675 477
<< mvpdiffc >>
rect -705 651 -699 657
rect -705 639 -699 645
rect -705 627 -699 633
rect -681 651 -675 657
rect -681 639 -675 645
rect -681 627 -675 633
<< psubdiff >>
rect -756 705 -660 708
rect -756 699 -753 705
rect -747 699 -741 705
rect -735 699 -729 705
rect -723 699 -717 705
rect -711 699 -705 705
rect -699 699 -693 705
rect -687 699 -681 705
rect -675 699 -669 705
rect -663 699 -660 705
rect -756 696 -660 699
rect -756 693 -744 696
rect -756 687 -753 693
rect -747 687 -744 693
rect -756 681 -744 687
rect -756 675 -753 681
rect -747 675 -744 681
rect -756 669 -744 675
rect -756 663 -753 669
rect -747 663 -744 669
rect -756 657 -744 663
rect -756 651 -753 657
rect -747 651 -744 657
rect -756 645 -744 651
rect -756 639 -753 645
rect -747 639 -744 645
rect -756 633 -744 639
rect -756 627 -753 633
rect -747 627 -744 633
rect -756 621 -744 627
rect -756 615 -753 621
rect -747 615 -744 621
rect -756 609 -744 615
rect -756 603 -753 609
rect -747 603 -744 609
rect -756 597 -744 603
rect -756 591 -753 597
rect -747 591 -744 597
rect -756 585 -744 591
rect -756 579 -753 585
rect -747 579 -744 585
rect -756 573 -744 579
rect -756 567 -753 573
rect -747 567 -744 573
rect -756 564 -744 567
rect -756 561 -660 564
rect -756 555 -753 561
rect -747 555 -741 561
rect -735 555 -729 561
rect -723 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -660 561
rect -756 552 -660 555
rect -756 549 -744 552
rect -756 543 -753 549
rect -747 543 -744 549
rect -756 537 -744 543
rect -756 531 -753 537
rect -747 531 -744 537
rect -756 525 -744 531
rect -756 519 -753 525
rect -747 519 -744 525
rect -756 513 -744 519
rect -756 507 -753 513
rect -747 507 -744 513
rect -756 501 -744 507
rect -756 495 -753 501
rect -747 495 -744 501
rect -756 489 -744 495
rect -756 483 -753 489
rect -747 483 -744 489
rect -756 477 -744 483
rect -756 471 -753 477
rect -747 471 -744 477
rect -756 465 -744 471
rect -756 459 -753 465
rect -747 459 -744 465
rect -756 453 -744 459
rect -756 447 -753 453
rect -747 447 -744 453
rect -756 441 -744 447
rect -756 435 -753 441
rect -747 435 -744 441
rect -756 429 -744 435
rect -756 423 -753 429
rect -747 423 -744 429
rect -756 417 -744 423
rect -756 411 -753 417
rect -747 411 -744 417
rect -756 408 -744 411
rect -756 405 -660 408
rect -756 399 -753 405
rect -747 399 -741 405
rect -735 399 -729 405
rect -723 399 -717 405
rect -711 399 -705 405
rect -699 399 -693 405
rect -687 399 -681 405
rect -675 399 -669 405
rect -663 399 -660 405
rect -756 396 -660 399
rect -756 393 -744 396
rect -756 387 -753 393
rect -747 387 -744 393
rect -756 381 -744 387
rect -756 375 -753 381
rect -747 375 -744 381
rect -756 357 -744 375
rect -756 351 -753 357
rect -747 351 -744 357
rect -756 345 -744 351
rect -756 339 -753 345
rect -747 339 -744 345
rect -756 333 -744 339
rect -756 327 -753 333
rect -747 327 -744 333
rect -756 309 -744 327
rect -756 303 -753 309
rect -747 303 -744 309
rect -756 297 -744 303
rect -756 291 -753 297
rect -747 291 -744 297
rect -756 288 -744 291
rect -756 285 -660 288
rect -756 279 -753 285
rect -747 279 -741 285
rect -735 279 -729 285
rect -723 279 -717 285
rect -711 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -669 285
rect -663 279 -660 285
rect -756 276 -660 279
rect -756 273 -744 276
rect -756 267 -753 273
rect -747 267 -744 273
rect -756 261 -744 267
rect -756 255 -753 261
rect -747 255 -744 261
rect -756 249 -744 255
rect -756 243 -753 249
rect -747 243 -744 249
rect -756 240 -744 243
rect -756 237 -660 240
rect -756 231 -753 237
rect -747 231 -741 237
rect -735 231 -729 237
rect -723 231 -717 237
rect -711 231 -705 237
rect -699 231 -693 237
rect -687 231 -681 237
rect -675 231 -669 237
rect -663 231 -660 237
rect -756 228 -660 231
rect -756 225 -744 228
rect -756 219 -753 225
rect -747 219 -744 225
rect -756 213 -744 219
rect -756 207 -753 213
rect -747 207 -744 213
rect -756 201 -744 207
rect -756 195 -753 201
rect -747 195 -744 201
rect -756 192 -744 195
rect -756 189 -660 192
rect -756 183 -753 189
rect -747 183 -741 189
rect -735 183 -729 189
rect -723 183 -717 189
rect -711 183 -705 189
rect -699 183 -693 189
rect -687 183 -681 189
rect -675 183 -669 189
rect -663 183 -660 189
rect -756 180 -660 183
rect -756 177 -744 180
rect -756 171 -753 177
rect -747 171 -744 177
rect -756 165 -744 171
rect -756 159 -753 165
rect -747 159 -744 165
rect -756 153 -744 159
rect -756 147 -753 153
rect -747 147 -744 153
rect -756 144 -744 147
rect -756 141 -660 144
rect -756 135 -753 141
rect -747 135 -741 141
rect -735 135 -729 141
rect -723 135 -717 141
rect -711 135 -705 141
rect -699 135 -693 141
rect -687 135 -681 141
rect -675 135 -669 141
rect -663 135 -660 141
rect -756 132 -660 135
rect -756 129 -744 132
rect -756 123 -753 129
rect -747 123 -744 129
rect -756 117 -744 123
rect -756 111 -753 117
rect -747 111 -744 117
rect -756 105 -744 111
rect -756 99 -753 105
rect -747 99 -744 105
rect -756 96 -744 99
rect -756 93 -660 96
rect -756 87 -753 93
rect -747 87 -741 93
rect -735 87 -729 93
rect -723 87 -717 93
rect -711 87 -705 93
rect -699 87 -693 93
rect -687 87 -681 93
rect -675 87 -669 93
rect -663 87 -660 93
rect -756 84 -660 87
rect -756 81 -744 84
rect -756 75 -753 81
rect -747 75 -744 81
rect -756 69 -744 75
rect -756 63 -753 69
rect -747 63 -744 69
rect -756 45 -744 63
rect -756 39 -753 45
rect -747 39 -744 45
rect -756 33 -744 39
rect -756 27 -753 33
rect -747 27 -744 33
rect -756 21 -744 27
rect -756 15 -753 21
rect -747 15 -744 21
rect -756 -3 -744 15
rect -756 -9 -753 -3
rect -747 -9 -744 -3
rect -756 -15 -744 -9
rect -756 -21 -753 -15
rect -747 -21 -744 -15
rect -756 -24 -744 -21
rect -756 -27 -660 -24
rect -756 -33 -753 -27
rect -747 -33 -741 -27
rect -735 -33 -729 -27
rect -723 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -39 -744 -36
rect -756 -45 -753 -39
rect -747 -45 -744 -39
rect -756 -51 -744 -45
rect -756 -57 -753 -51
rect -747 -57 -744 -51
rect -756 -63 -744 -57
rect -756 -69 -753 -63
rect -747 -69 -744 -63
rect -756 -75 -744 -69
rect -756 -81 -753 -75
rect -747 -81 -744 -75
rect -756 -87 -744 -81
rect -756 -93 -753 -87
rect -747 -93 -744 -87
rect -756 -99 -744 -93
rect -756 -105 -753 -99
rect -747 -105 -744 -99
rect -756 -111 -744 -105
rect -756 -117 -753 -111
rect -747 -117 -744 -111
rect -756 -120 -744 -117
rect -756 -123 -660 -120
rect -756 -129 -753 -123
rect -747 -129 -741 -123
rect -735 -129 -729 -123
rect -723 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -660 -123
rect -756 -132 -660 -129
<< nsubdiff >>
rect -732 537 -672 540
rect -732 531 -729 537
rect -723 531 -717 537
rect -711 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -672 537
rect -732 528 -672 531
rect -732 525 -720 528
rect -732 519 -729 525
rect -723 519 -720 525
rect -732 513 -720 519
rect -732 507 -729 513
rect -723 507 -720 513
rect -732 501 -720 507
rect -732 495 -729 501
rect -723 495 -720 501
rect -732 489 -720 495
rect -732 483 -729 489
rect -723 483 -720 489
rect -732 477 -720 483
rect -732 471 -729 477
rect -723 471 -720 477
rect -732 465 -720 471
rect -732 459 -729 465
rect -723 459 -720 465
rect -732 453 -720 459
rect -732 447 -729 453
rect -723 447 -720 453
rect -732 441 -720 447
rect -732 435 -729 441
rect -723 435 -720 441
rect -732 432 -720 435
rect -732 429 -672 432
rect -732 423 -729 429
rect -723 423 -717 429
rect -711 423 -705 429
rect -699 423 -693 429
rect -687 423 -681 429
rect -675 423 -672 429
rect -732 420 -672 423
<< mvnsubdiff >>
rect -732 681 -672 684
rect -732 675 -729 681
rect -723 675 -717 681
rect -711 675 -705 681
rect -699 675 -693 681
rect -687 675 -681 681
rect -675 675 -672 681
rect -732 672 -672 675
rect -732 669 -720 672
rect -732 663 -729 669
rect -723 663 -720 669
rect -732 657 -720 663
rect -732 651 -729 657
rect -723 651 -720 657
rect -732 645 -720 651
rect -732 639 -729 645
rect -723 639 -720 645
rect -732 633 -720 639
rect -732 627 -729 633
rect -723 627 -720 633
rect -732 621 -720 627
rect -732 615 -729 621
rect -723 615 -720 621
rect -732 609 -720 615
rect -732 603 -729 609
rect -723 603 -720 609
rect -732 597 -720 603
rect -732 591 -729 597
rect -723 591 -720 597
rect -732 588 -720 591
rect -732 585 -672 588
rect -732 579 -729 585
rect -723 579 -717 585
rect -711 579 -705 585
rect -699 579 -693 585
rect -687 579 -681 585
rect -675 579 -672 585
rect -732 576 -672 579
<< psubdiffcont >>
rect -753 699 -747 705
rect -741 699 -735 705
rect -729 699 -723 705
rect -717 699 -711 705
rect -705 699 -699 705
rect -693 699 -687 705
rect -681 699 -675 705
rect -669 699 -663 705
rect -753 687 -747 693
rect -753 675 -747 681
rect -753 663 -747 669
rect -753 651 -747 657
rect -753 639 -747 645
rect -753 627 -747 633
rect -753 615 -747 621
rect -753 603 -747 609
rect -753 591 -747 597
rect -753 579 -747 585
rect -753 567 -747 573
rect -753 555 -747 561
rect -741 555 -735 561
rect -729 555 -723 561
rect -717 555 -711 561
rect -705 555 -699 561
rect -693 555 -687 561
rect -681 555 -675 561
rect -669 555 -663 561
rect -753 543 -747 549
rect -753 531 -747 537
rect -753 519 -747 525
rect -753 507 -747 513
rect -753 495 -747 501
rect -753 483 -747 489
rect -753 471 -747 477
rect -753 459 -747 465
rect -753 447 -747 453
rect -753 435 -747 441
rect -753 423 -747 429
rect -753 411 -747 417
rect -753 399 -747 405
rect -741 399 -735 405
rect -729 399 -723 405
rect -717 399 -711 405
rect -705 399 -699 405
rect -693 399 -687 405
rect -681 399 -675 405
rect -669 399 -663 405
rect -753 387 -747 393
rect -753 375 -747 381
rect -753 351 -747 357
rect -753 339 -747 345
rect -753 327 -747 333
rect -753 303 -747 309
rect -753 291 -747 297
rect -753 279 -747 285
rect -741 279 -735 285
rect -729 279 -723 285
rect -717 279 -711 285
rect -705 279 -699 285
rect -693 279 -687 285
rect -681 279 -675 285
rect -669 279 -663 285
rect -753 267 -747 273
rect -753 255 -747 261
rect -753 243 -747 249
rect -753 231 -747 237
rect -741 231 -735 237
rect -729 231 -723 237
rect -717 231 -711 237
rect -705 231 -699 237
rect -693 231 -687 237
rect -681 231 -675 237
rect -669 231 -663 237
rect -753 219 -747 225
rect -753 207 -747 213
rect -753 195 -747 201
rect -753 183 -747 189
rect -741 183 -735 189
rect -729 183 -723 189
rect -717 183 -711 189
rect -705 183 -699 189
rect -693 183 -687 189
rect -681 183 -675 189
rect -669 183 -663 189
rect -753 171 -747 177
rect -753 159 -747 165
rect -753 147 -747 153
rect -753 135 -747 141
rect -741 135 -735 141
rect -729 135 -723 141
rect -717 135 -711 141
rect -705 135 -699 141
rect -693 135 -687 141
rect -681 135 -675 141
rect -669 135 -663 141
rect -753 123 -747 129
rect -753 111 -747 117
rect -753 99 -747 105
rect -753 87 -747 93
rect -741 87 -735 93
rect -729 87 -723 93
rect -717 87 -711 93
rect -705 87 -699 93
rect -693 87 -687 93
rect -681 87 -675 93
rect -669 87 -663 93
rect -753 75 -747 81
rect -753 63 -747 69
rect -753 39 -747 45
rect -753 27 -747 33
rect -753 15 -747 21
rect -753 -9 -747 -3
rect -753 -21 -747 -15
rect -753 -33 -747 -27
rect -741 -33 -735 -27
rect -729 -33 -723 -27
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -753 -45 -747 -39
rect -753 -57 -747 -51
rect -753 -69 -747 -63
rect -753 -81 -747 -75
rect -753 -93 -747 -87
rect -753 -105 -747 -99
rect -753 -117 -747 -111
rect -753 -129 -747 -123
rect -741 -129 -735 -123
rect -729 -129 -723 -123
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
<< nsubdiffcont >>
rect -729 531 -723 537
rect -717 531 -711 537
rect -705 531 -699 537
rect -693 531 -687 537
rect -681 531 -675 537
rect -729 519 -723 525
rect -729 507 -723 513
rect -729 495 -723 501
rect -729 483 -723 489
rect -729 471 -723 477
rect -729 459 -723 465
rect -729 447 -723 453
rect -729 435 -723 441
rect -729 423 -723 429
rect -717 423 -711 429
rect -705 423 -699 429
rect -693 423 -687 429
rect -681 423 -675 429
<< mvnsubdiffcont >>
rect -729 675 -723 681
rect -717 675 -711 681
rect -705 675 -699 681
rect -693 675 -687 681
rect -681 675 -675 681
rect -729 663 -723 669
rect -729 651 -723 657
rect -729 639 -723 645
rect -729 627 -723 633
rect -729 615 -723 621
rect -729 603 -723 609
rect -729 591 -723 597
rect -729 579 -723 585
rect -717 579 -711 585
rect -705 579 -699 585
rect -693 579 -687 585
rect -681 579 -675 585
<< polysilicon >>
rect -696 660 -684 666
rect -696 609 -684 624
rect -696 603 -693 609
rect -687 603 -684 609
rect -696 600 -684 603
rect -696 498 -684 504
rect -696 453 -684 468
rect -696 447 -693 453
rect -687 447 -684 453
rect -696 444 -684 447
rect -696 -51 -684 -48
rect -696 -57 -693 -51
rect -687 -57 -684 -51
rect -696 -72 -684 -57
rect -696 -114 -684 -108
<< polycontact >>
rect -693 603 -687 609
rect -693 447 -687 453
rect -693 -57 -687 -51
<< metal1 >>
rect -756 705 -660 708
rect -756 699 -753 705
rect -747 699 -741 705
rect -735 699 -729 705
rect -723 699 -717 705
rect -711 699 -705 705
rect -699 699 -693 705
rect -687 699 -681 705
rect -675 699 -669 705
rect -663 699 -660 705
rect -756 696 -660 699
rect -756 693 -744 696
rect -756 687 -753 693
rect -747 687 -744 693
rect -756 681 -744 687
rect -756 675 -753 681
rect -747 675 -744 681
rect -756 669 -744 675
rect -756 663 -753 669
rect -747 663 -744 669
rect -756 657 -744 663
rect -756 651 -753 657
rect -747 651 -744 657
rect -756 645 -744 651
rect -756 639 -753 645
rect -747 639 -744 645
rect -756 633 -744 639
rect -756 627 -753 633
rect -747 627 -744 633
rect -756 621 -744 627
rect -756 615 -753 621
rect -747 615 -744 621
rect -756 609 -744 615
rect -756 603 -753 609
rect -747 603 -744 609
rect -756 597 -744 603
rect -756 591 -753 597
rect -747 591 -744 597
rect -756 585 -744 591
rect -756 579 -753 585
rect -747 579 -744 585
rect -756 573 -744 579
rect -732 681 -660 684
rect -732 675 -729 681
rect -723 675 -717 681
rect -711 675 -705 681
rect -699 675 -693 681
rect -687 675 -681 681
rect -675 675 -660 681
rect -732 672 -660 675
rect -732 669 -720 672
rect -732 663 -729 669
rect -723 663 -720 669
rect -732 657 -720 663
rect -732 651 -729 657
rect -723 651 -720 657
rect -732 645 -720 651
rect -732 639 -729 645
rect -723 639 -720 645
rect -732 633 -720 639
rect -732 627 -729 633
rect -723 627 -720 633
rect -732 621 -720 627
rect -732 615 -729 621
rect -723 615 -720 621
rect -732 609 -720 615
rect -732 603 -729 609
rect -723 603 -720 609
rect -732 597 -720 603
rect -708 657 -696 660
rect -708 651 -705 657
rect -699 651 -696 657
rect -708 645 -696 651
rect -708 639 -705 645
rect -699 639 -696 645
rect -708 633 -696 639
rect -708 627 -705 633
rect -699 627 -696 633
rect -708 612 -696 627
rect -684 657 -672 660
rect -684 651 -681 657
rect -675 651 -672 657
rect -684 645 -672 651
rect -684 639 -681 645
rect -675 639 -672 645
rect -684 633 -672 639
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 624 -672 627
rect -708 609 -684 612
rect -708 603 -693 609
rect -687 603 -684 609
rect -708 600 -684 603
rect -732 591 -729 597
rect -723 591 -720 597
rect -732 588 -720 591
rect -732 585 -660 588
rect -732 579 -729 585
rect -723 579 -717 585
rect -711 579 -705 585
rect -699 579 -693 585
rect -687 579 -681 585
rect -675 579 -660 585
rect -732 576 -660 579
rect -756 567 -753 573
rect -747 567 -744 573
rect -756 564 -744 567
rect -756 561 -660 564
rect -756 555 -753 561
rect -747 555 -741 561
rect -735 555 -729 561
rect -723 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -660 561
rect -756 552 -660 555
rect -756 549 -744 552
rect -756 543 -753 549
rect -747 543 -744 549
rect -756 537 -744 543
rect -756 531 -753 537
rect -747 531 -744 537
rect -756 525 -744 531
rect -756 519 -753 525
rect -747 519 -744 525
rect -756 513 -744 519
rect -756 507 -753 513
rect -747 507 -744 513
rect -756 501 -744 507
rect -756 495 -753 501
rect -747 495 -744 501
rect -756 489 -744 495
rect -756 483 -753 489
rect -747 483 -744 489
rect -756 477 -744 483
rect -756 471 -753 477
rect -747 471 -744 477
rect -756 465 -744 471
rect -756 459 -753 465
rect -747 459 -744 465
rect -756 453 -744 459
rect -756 447 -753 453
rect -747 447 -744 453
rect -756 441 -744 447
rect -756 435 -753 441
rect -747 435 -744 441
rect -756 429 -744 435
rect -756 423 -753 429
rect -747 423 -744 429
rect -756 417 -744 423
rect -732 537 -672 540
rect -732 531 -729 537
rect -723 531 -717 537
rect -711 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -672 537
rect -732 528 -672 531
rect -732 525 -720 528
rect -732 519 -729 525
rect -723 519 -720 525
rect -732 513 -720 519
rect -732 507 -729 513
rect -723 507 -720 513
rect -732 501 -720 507
rect -732 495 -729 501
rect -723 495 -720 501
rect -732 489 -720 495
rect -732 483 -729 489
rect -723 483 -720 489
rect -732 477 -720 483
rect -732 471 -729 477
rect -723 471 -720 477
rect -732 465 -720 471
rect -732 459 -729 465
rect -723 459 -720 465
rect -732 453 -720 459
rect -732 447 -729 453
rect -723 447 -720 453
rect -732 441 -720 447
rect -708 489 -696 498
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 477 -696 483
rect -708 471 -705 477
rect -699 471 -696 477
rect -708 456 -696 471
rect -684 489 -672 498
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 477 -672 483
rect -684 471 -681 477
rect -675 471 -672 477
rect -684 468 -672 471
rect -708 453 -684 456
rect -708 447 -693 453
rect -687 447 -684 453
rect -708 444 -684 447
rect -732 435 -729 441
rect -723 435 -720 441
rect -732 432 -720 435
rect -732 429 -660 432
rect -732 423 -729 429
rect -723 423 -717 429
rect -711 423 -705 429
rect -699 423 -693 429
rect -687 423 -681 429
rect -675 423 -660 429
rect -732 420 -660 423
rect -756 411 -753 417
rect -747 411 -744 417
rect -756 408 -744 411
rect -756 405 -660 408
rect -756 399 -753 405
rect -747 399 -741 405
rect -735 399 -729 405
rect -723 399 -717 405
rect -711 399 -705 405
rect -699 399 -693 405
rect -687 399 -681 405
rect -675 399 -669 405
rect -663 399 -660 405
rect -756 396 -660 399
rect -756 393 -744 396
rect -756 387 -753 393
rect -747 387 -744 393
rect -756 381 -744 387
rect -756 375 -753 381
rect -747 375 -744 381
rect -756 357 -744 375
rect -756 351 -753 357
rect -747 351 -744 357
rect -756 345 -744 351
rect -756 339 -753 345
rect -747 339 -744 345
rect -756 333 -744 339
rect -756 327 -753 333
rect -747 327 -744 333
rect -756 309 -744 327
rect -756 303 -753 309
rect -747 303 -744 309
rect -756 297 -744 303
rect -756 291 -753 297
rect -747 291 -744 297
rect -756 288 -744 291
rect -756 285 -660 288
rect -756 279 -753 285
rect -747 279 -741 285
rect -735 279 -729 285
rect -723 279 -717 285
rect -711 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -669 285
rect -663 279 -660 285
rect -756 276 -660 279
rect -756 273 -744 276
rect -756 267 -753 273
rect -747 267 -744 273
rect -756 261 -744 267
rect -756 255 -753 261
rect -747 255 -744 261
rect -756 249 -744 255
rect -756 243 -753 249
rect -747 243 -744 249
rect -756 240 -744 243
rect -756 237 -660 240
rect -756 231 -753 237
rect -747 231 -741 237
rect -735 231 -729 237
rect -723 231 -717 237
rect -711 231 -705 237
rect -699 231 -693 237
rect -687 231 -681 237
rect -675 231 -669 237
rect -663 231 -660 237
rect -756 228 -660 231
rect -756 225 -744 228
rect -756 219 -753 225
rect -747 219 -744 225
rect -756 213 -744 219
rect -756 207 -753 213
rect -747 207 -744 213
rect -756 201 -744 207
rect -756 195 -753 201
rect -747 195 -744 201
rect -756 192 -744 195
rect -756 189 -660 192
rect -756 183 -753 189
rect -747 183 -741 189
rect -735 183 -729 189
rect -723 183 -717 189
rect -711 183 -705 189
rect -699 183 -693 189
rect -687 183 -681 189
rect -675 183 -669 189
rect -663 183 -660 189
rect -756 180 -660 183
rect -756 177 -744 180
rect -756 171 -753 177
rect -747 171 -744 177
rect -756 165 -744 171
rect -756 159 -753 165
rect -747 159 -744 165
rect -756 153 -744 159
rect -756 147 -753 153
rect -747 147 -744 153
rect -756 144 -744 147
rect -756 141 -660 144
rect -756 135 -753 141
rect -747 135 -741 141
rect -735 135 -729 141
rect -723 135 -717 141
rect -711 135 -705 141
rect -699 135 -693 141
rect -687 135 -681 141
rect -675 135 -669 141
rect -663 135 -660 141
rect -756 132 -660 135
rect -756 129 -744 132
rect -756 123 -753 129
rect -747 123 -744 129
rect -756 117 -744 123
rect -756 111 -753 117
rect -747 111 -744 117
rect -756 105 -744 111
rect -756 99 -753 105
rect -747 99 -744 105
rect -756 96 -744 99
rect -756 93 -660 96
rect -756 87 -753 93
rect -747 87 -741 93
rect -735 87 -729 93
rect -723 87 -717 93
rect -711 87 -705 93
rect -699 87 -693 93
rect -687 87 -681 93
rect -675 87 -669 93
rect -663 87 -660 93
rect -756 84 -660 87
rect -756 81 -744 84
rect -756 75 -753 81
rect -747 75 -744 81
rect -756 69 -744 75
rect -756 63 -753 69
rect -747 63 -744 69
rect -756 45 -744 63
rect -756 39 -753 45
rect -747 39 -744 45
rect -756 33 -744 39
rect -756 27 -753 33
rect -747 27 -744 33
rect -756 21 -744 27
rect -756 15 -753 21
rect -747 15 -744 21
rect -756 -3 -744 15
rect -756 -9 -753 -3
rect -747 -9 -744 -3
rect -756 -15 -744 -9
rect -756 -21 -753 -15
rect -747 -21 -744 -15
rect -756 -24 -744 -21
rect -756 -27 -660 -24
rect -756 -33 -753 -27
rect -747 -33 -741 -27
rect -735 -33 -729 -27
rect -723 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -39 -744 -36
rect -756 -45 -753 -39
rect -747 -45 -744 -39
rect -756 -51 -744 -45
rect -756 -57 -753 -51
rect -747 -57 -744 -51
rect -756 -63 -744 -57
rect -756 -69 -753 -63
rect -747 -69 -744 -63
rect -756 -75 -744 -69
rect -756 -81 -753 -75
rect -747 -81 -744 -75
rect -756 -87 -744 -81
rect -756 -93 -753 -87
rect -747 -93 -744 -87
rect -756 -99 -744 -93
rect -756 -105 -753 -99
rect -747 -105 -744 -99
rect -756 -111 -744 -105
rect -708 -51 -684 -48
rect -708 -57 -693 -51
rect -687 -57 -684 -51
rect -708 -60 -684 -57
rect -708 -75 -696 -60
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -756 -117 -753 -111
rect -747 -117 -744 -111
rect -756 -120 -744 -117
rect -756 -123 -660 -120
rect -756 -129 -753 -123
rect -747 -129 -741 -123
rect -735 -129 -729 -123
rect -723 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -660 -123
rect -756 -132 -660 -129
<< via1 >>
rect -681 675 -675 681
rect -681 651 -675 657
rect -681 639 -675 645
rect -681 627 -675 633
rect -681 483 -675 489
rect -681 471 -675 477
rect -729 423 -723 429
rect -681 399 -675 405
rect -681 279 -675 285
rect -681 231 -675 237
rect -681 183 -675 189
rect -681 135 -675 141
rect -681 87 -675 93
rect -681 -33 -675 -27
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -681 -129 -675 -123
<< metal2 >>
rect -684 681 -672 684
rect -684 675 -681 681
rect -675 675 -672 681
rect -684 657 -672 675
rect -684 651 -681 657
rect -675 651 -672 657
rect -684 645 -672 651
rect -684 639 -681 645
rect -675 639 -672 645
rect -684 633 -672 639
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 624 -672 627
rect -708 585 -696 588
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 537 -696 579
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 528 -696 531
rect -684 537 -672 540
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 489 -672 531
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 477 -672 483
rect -684 471 -681 477
rect -675 471 -672 477
rect -684 468 -672 471
rect -732 429 -720 432
rect -732 423 -729 429
rect -723 423 -720 429
rect -732 420 -720 423
rect -684 405 -672 408
rect -684 399 -681 405
rect -675 399 -672 405
rect -684 285 -672 399
rect -684 279 -681 285
rect -675 279 -672 285
rect -684 237 -672 279
rect -684 231 -681 237
rect -675 231 -672 237
rect -684 189 -672 231
rect -684 183 -681 189
rect -675 183 -672 189
rect -684 141 -672 183
rect -684 135 -681 141
rect -675 135 -672 141
rect -684 93 -672 135
rect -684 87 -681 93
rect -675 87 -672 93
rect -684 -27 -672 87
rect -684 -33 -681 -27
rect -675 -33 -672 -27
rect -684 -75 -672 -33
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -123 -672 -105
rect -684 -129 -681 -123
rect -675 -129 -672 -123
rect -684 -132 -672 -129
<< via2 >>
rect -681 675 -675 681
rect -681 651 -675 657
rect -681 639 -675 645
rect -681 627 -675 633
rect -705 579 -699 585
rect -705 531 -699 537
rect -681 531 -675 537
rect -729 423 -723 429
rect -681 399 -675 405
rect -681 279 -675 285
rect -681 231 -675 237
rect -681 183 -675 189
rect -681 135 -675 141
rect -681 87 -675 93
rect -681 -33 -675 -27
rect -681 -129 -675 -123
<< metal3 >>
rect -756 681 -660 684
rect -756 675 -681 681
rect -675 675 -660 681
rect -756 657 -660 675
rect -756 651 -681 657
rect -675 651 -660 657
rect -756 645 -660 651
rect -756 639 -681 645
rect -675 639 -660 645
rect -756 633 -660 639
rect -756 627 -681 633
rect -675 627 -660 633
rect -756 624 -660 627
rect -756 585 -660 588
rect -756 579 -705 585
rect -699 579 -660 585
rect -756 570 -660 579
rect -756 552 -660 564
rect -756 537 -660 546
rect -756 531 -705 537
rect -699 531 -681 537
rect -675 531 -660 537
rect -756 528 -660 531
rect -756 429 -660 432
rect -756 423 -729 429
rect -723 423 -660 429
rect -756 420 -660 423
rect -756 405 -660 408
rect -756 399 -681 405
rect -675 399 -660 405
rect -756 396 -660 399
rect -756 354 -660 384
rect -756 336 -660 348
rect -756 300 -660 330
rect -756 285 -660 288
rect -756 279 -681 285
rect -675 279 -660 285
rect -756 276 -660 279
rect -756 252 -660 264
rect -756 237 -660 240
rect -756 231 -681 237
rect -675 231 -660 237
rect -756 228 -660 231
rect -756 204 -660 216
rect -756 189 -660 192
rect -756 183 -681 189
rect -675 183 -660 189
rect -756 180 -660 183
rect -756 156 -660 168
rect -756 141 -660 144
rect -756 135 -681 141
rect -675 135 -660 141
rect -756 132 -660 135
rect -756 108 -660 120
rect -756 93 -660 96
rect -756 87 -681 93
rect -675 87 -660 93
rect -756 84 -660 87
rect -756 42 -660 72
rect -756 24 -660 36
rect -756 -12 -660 18
rect -756 -27 -660 -24
rect -756 -33 -681 -27
rect -675 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -123 -660 -72
rect -756 -129 -681 -123
rect -675 -129 -660 -123
rect -756 -132 -660 -129
<< labels >>
rlabel metal3 -756 -132 -660 -72 0 gnd
port 9 nsew
rlabel metal1 -708 -60 -696 -48 0 lo
rlabel metal3 -756 -12 -660 0 0 om
port 13 nsew
rlabel metal3 -756 24 -660 36 0 xp
port 12 nsew
rlabel metal3 -756 108 -660 120 0 ip
port 7 nsew
rlabel metal3 -756 60 -660 72 0 om
port 13 nsew
rlabel metal3 -756 252 -660 264 0 im
port 6 nsew
rlabel metal3 -756 336 -660 348 0 xm
port 10 nsew
rlabel metal3 -756 372 -660 384 0 op
port 11 nsew
rlabel metal1 -708 444 -696 456 0 hi
rlabel metal1 -708 600 -696 612 1 hih
rlabel metal3 -756 576 -660 588 0 vreg
port 4 nsew
rlabel metal3 -756 420 -660 432 0 bp
port 3 nsew
rlabel metal3 -756 552 -660 564 0 gp
port 2 nsew
rlabel metal3 -756 624 -660 684 0 vdd
port 1 nsew
rlabel metal3 -756 300 -660 312 0 op
port 11 nsew
rlabel metal3 -756 204 -660 216 0 x
port 14 nsew
rlabel metal3 -756 156 -660 168 0 y
port 15 nsew
<< end >>
