magic
tech gf180mcuC
timestamp 1665298770
<< via2 >>
rect -408 228 -396 252
rect -48 228 -36 252
rect 192 228 204 252
rect 312 228 324 252
rect 552 228 564 252
rect 912 228 924 252
rect 1032 228 1044 252
rect 1392 228 1404 252
rect 1632 228 1644 252
rect 1752 228 1764 252
rect 1992 228 2004 252
rect 2352 228 2364 252
rect -648 204 -636 216
rect -528 204 -516 216
rect 2472 204 2484 216
rect 2592 204 2604 216
rect -408 168 -396 192
rect -48 168 -36 192
rect 192 168 204 192
rect 312 168 324 192
rect 552 168 564 192
rect 912 168 924 192
rect 1032 168 1044 192
rect 1392 168 1404 192
rect 1632 168 1644 192
rect 1752 168 1764 192
rect 1992 168 2004 192
rect 2352 168 2364 192
rect -288 12 -276 36
rect -168 12 -156 36
rect 72 12 84 36
rect 432 12 444 36
rect 672 12 684 36
rect 792 12 804 36
rect 1152 12 1164 36
rect 1272 12 1284 36
rect 1512 12 1524 36
rect 1872 12 1884 36
rect 2112 12 2124 36
rect 2232 12 2244 36
rect -888 -12 -876 0
rect -768 -12 -756 0
rect 2712 -12 2724 0
rect 2832 -12 2844 0
rect -288 -48 -276 -24
rect -168 -48 -156 -24
rect 72 -48 84 -24
rect 432 -48 444 -24
rect 672 -48 684 -24
rect 792 -48 804 -24
rect 1152 -48 1164 -24
rect 1272 -48 1284 -24
rect 1512 -48 1524 -24
rect 1872 -48 1884 -24
rect 2112 -48 2124 -24
rect 2232 -48 2244 -24
<< mimcap >>
rect -1008 792 2976 804
rect -1008 780 -996 792
rect -984 780 -972 792
rect -960 780 -948 792
rect -936 780 -924 792
rect -912 780 -900 792
rect -888 780 -876 792
rect -864 780 -852 792
rect -840 780 -828 792
rect -816 780 -804 792
rect -792 780 -780 792
rect -768 780 -756 792
rect -744 780 -732 792
rect -720 780 -708 792
rect -696 780 -684 792
rect -672 780 -660 792
rect -648 780 -636 792
rect -624 780 -612 792
rect -600 780 -588 792
rect -576 780 -564 792
rect -552 780 -540 792
rect -528 780 -516 792
rect -504 780 -492 792
rect -480 780 -468 792
rect -456 780 -444 792
rect -432 780 -420 792
rect -408 780 -396 792
rect -384 780 -372 792
rect -360 780 -348 792
rect -336 780 -324 792
rect -312 780 -300 792
rect -288 780 -276 792
rect -264 780 -252 792
rect -240 780 -228 792
rect -216 780 -204 792
rect -192 780 -180 792
rect -168 780 -156 792
rect -144 780 -132 792
rect -120 780 -108 792
rect -96 780 -84 792
rect -72 780 -60 792
rect -48 780 -36 792
rect -24 780 -12 792
rect 0 780 12 792
rect 24 780 36 792
rect 48 780 60 792
rect 72 780 84 792
rect 96 780 108 792
rect 120 780 132 792
rect 144 780 156 792
rect 168 780 180 792
rect 192 780 204 792
rect 216 780 228 792
rect 240 780 252 792
rect 264 780 276 792
rect 288 780 300 792
rect 312 780 324 792
rect 336 780 348 792
rect 360 780 372 792
rect 384 780 396 792
rect 408 780 420 792
rect 432 780 444 792
rect 456 780 468 792
rect 480 780 492 792
rect 504 780 516 792
rect 528 780 540 792
rect 552 780 564 792
rect 576 780 588 792
rect 600 780 612 792
rect 624 780 636 792
rect 648 780 660 792
rect 672 780 684 792
rect 696 780 708 792
rect 720 780 732 792
rect 744 780 756 792
rect 768 780 780 792
rect 792 780 804 792
rect 816 780 828 792
rect 840 780 852 792
rect 864 780 876 792
rect 888 780 900 792
rect 912 780 924 792
rect 936 780 948 792
rect 960 780 972 792
rect 984 780 996 792
rect 1008 780 1020 792
rect 1032 780 1044 792
rect 1056 780 1068 792
rect 1080 780 1092 792
rect 1104 780 1116 792
rect 1128 780 1140 792
rect 1152 780 1164 792
rect 1176 780 1188 792
rect 1200 780 1212 792
rect 1224 780 1236 792
rect 1248 780 1260 792
rect 1272 780 1284 792
rect 1296 780 1308 792
rect 1320 780 1332 792
rect 1344 780 1356 792
rect 1368 780 1380 792
rect 1392 780 1404 792
rect 1416 780 1428 792
rect 1440 780 1452 792
rect 1464 780 1476 792
rect 1488 780 1500 792
rect 1512 780 1524 792
rect 1536 780 1548 792
rect 1560 780 1572 792
rect 1584 780 1596 792
rect 1608 780 1620 792
rect 1632 780 1644 792
rect 1656 780 1668 792
rect 1680 780 1692 792
rect 1704 780 1716 792
rect 1728 780 1740 792
rect 1752 780 1764 792
rect 1776 780 1788 792
rect 1800 780 1812 792
rect 1824 780 1836 792
rect 1848 780 1860 792
rect 1872 780 1884 792
rect 1896 780 1908 792
rect 1920 780 1932 792
rect 1944 780 1956 792
rect 1968 780 1980 792
rect 1992 780 2004 792
rect 2016 780 2028 792
rect 2040 780 2052 792
rect 2064 780 2076 792
rect 2088 780 2100 792
rect 2112 780 2124 792
rect 2136 780 2148 792
rect 2160 780 2172 792
rect 2184 780 2196 792
rect 2208 780 2220 792
rect 2232 780 2244 792
rect 2256 780 2268 792
rect 2280 780 2292 792
rect 2304 780 2316 792
rect 2328 780 2340 792
rect 2352 780 2364 792
rect 2376 780 2388 792
rect 2400 780 2412 792
rect 2424 780 2436 792
rect 2448 780 2460 792
rect 2472 780 2484 792
rect 2496 780 2508 792
rect 2520 780 2532 792
rect 2544 780 2556 792
rect 2568 780 2580 792
rect 2592 780 2604 792
rect 2616 780 2628 792
rect 2640 780 2652 792
rect 2664 780 2676 792
rect 2688 780 2700 792
rect 2712 780 2724 792
rect 2736 780 2748 792
rect 2760 780 2772 792
rect 2784 780 2796 792
rect 2808 780 2820 792
rect 2832 780 2844 792
rect 2856 780 2868 792
rect 2880 780 2892 792
rect 2904 780 2916 792
rect 2928 780 2940 792
rect 2952 780 2976 792
rect -1008 756 2976 780
rect -1008 744 -996 756
rect -984 744 -972 756
rect -960 744 -948 756
rect -936 744 -924 756
rect -912 744 -900 756
rect -888 744 -876 756
rect -864 744 -852 756
rect -840 744 -828 756
rect -816 744 -804 756
rect -792 744 -780 756
rect -768 744 -756 756
rect -744 744 -732 756
rect -720 744 -708 756
rect -696 744 -684 756
rect -672 744 -660 756
rect -648 744 -636 756
rect -624 744 -612 756
rect -600 744 -588 756
rect -576 744 -564 756
rect -552 744 -540 756
rect -528 744 -516 756
rect -504 744 -492 756
rect -480 744 -468 756
rect -456 744 -444 756
rect -432 744 -420 756
rect -408 744 -396 756
rect -384 744 -372 756
rect -360 744 -348 756
rect -336 744 -324 756
rect -312 744 -300 756
rect -288 744 -276 756
rect -264 744 -252 756
rect -240 744 -228 756
rect -216 744 -204 756
rect -192 744 -180 756
rect -168 744 -156 756
rect -144 744 -132 756
rect -120 744 -108 756
rect -96 744 -84 756
rect -72 744 -60 756
rect -48 744 -36 756
rect -24 744 -12 756
rect 0 744 12 756
rect 24 744 36 756
rect 48 744 60 756
rect 72 744 84 756
rect 96 744 108 756
rect 120 744 132 756
rect 144 744 156 756
rect 168 744 180 756
rect 192 744 204 756
rect 216 744 228 756
rect 240 744 252 756
rect 264 744 276 756
rect 288 744 300 756
rect 312 744 324 756
rect 336 744 348 756
rect 360 744 372 756
rect 384 744 396 756
rect 408 744 420 756
rect 432 744 444 756
rect 456 744 468 756
rect 480 744 492 756
rect 504 744 516 756
rect 528 744 540 756
rect 552 744 564 756
rect 576 744 588 756
rect 600 744 612 756
rect 624 744 636 756
rect 648 744 660 756
rect 672 744 684 756
rect 696 744 708 756
rect 720 744 732 756
rect 744 744 756 756
rect 768 744 780 756
rect 792 744 804 756
rect 816 744 828 756
rect 840 744 852 756
rect 864 744 876 756
rect 888 744 900 756
rect 912 744 924 756
rect 936 744 948 756
rect 960 744 972 756
rect 984 744 996 756
rect 1008 744 1020 756
rect 1032 744 1044 756
rect 1056 744 1068 756
rect 1080 744 1092 756
rect 1104 744 1116 756
rect 1128 744 1140 756
rect 1152 744 1164 756
rect 1176 744 1188 756
rect 1200 744 1212 756
rect 1224 744 1236 756
rect 1248 744 1260 756
rect 1272 744 1284 756
rect 1296 744 1308 756
rect 1320 744 1332 756
rect 1344 744 1356 756
rect 1368 744 1380 756
rect 1392 744 1404 756
rect 1416 744 1428 756
rect 1440 744 1452 756
rect 1464 744 1476 756
rect 1488 744 1500 756
rect 1512 744 1524 756
rect 1536 744 1548 756
rect 1560 744 1572 756
rect 1584 744 1596 756
rect 1608 744 1620 756
rect 1632 744 1644 756
rect 1656 744 1668 756
rect 1680 744 1692 756
rect 1704 744 1716 756
rect 1728 744 1740 756
rect 1752 744 1764 756
rect 1776 744 1788 756
rect 1800 744 1812 756
rect 1824 744 1836 756
rect 1848 744 1860 756
rect 1872 744 1884 756
rect 1896 744 1908 756
rect 1920 744 1932 756
rect 1944 744 1956 756
rect 1968 744 1980 756
rect 1992 744 2004 756
rect 2016 744 2028 756
rect 2040 744 2052 756
rect 2064 744 2076 756
rect 2088 744 2100 756
rect 2112 744 2124 756
rect 2136 744 2148 756
rect 2160 744 2172 756
rect 2184 744 2196 756
rect 2208 744 2220 756
rect 2232 744 2244 756
rect 2256 744 2268 756
rect 2280 744 2292 756
rect 2304 744 2316 756
rect 2328 744 2340 756
rect 2352 744 2364 756
rect 2376 744 2388 756
rect 2400 744 2412 756
rect 2424 744 2436 756
rect 2448 744 2460 756
rect 2472 744 2484 756
rect 2496 744 2508 756
rect 2520 744 2532 756
rect 2544 744 2556 756
rect 2568 744 2580 756
rect 2592 744 2604 756
rect 2616 744 2628 756
rect 2640 744 2652 756
rect 2664 744 2676 756
rect 2688 744 2700 756
rect 2712 744 2724 756
rect 2736 744 2748 756
rect 2760 744 2772 756
rect 2784 744 2796 756
rect 2808 744 2820 756
rect 2832 744 2844 756
rect 2856 744 2868 756
rect 2880 744 2892 756
rect 2904 744 2916 756
rect 2928 744 2940 756
rect 2952 744 2976 756
rect -1008 720 2976 744
rect -1008 708 -996 720
rect -984 708 -972 720
rect -960 708 -948 720
rect -936 708 -924 720
rect -912 708 -900 720
rect -888 708 -876 720
rect -864 708 -852 720
rect -840 708 -828 720
rect -816 708 -804 720
rect -792 708 -780 720
rect -768 708 -756 720
rect -744 708 -732 720
rect -720 708 -708 720
rect -696 708 -684 720
rect -672 708 -660 720
rect -648 708 -636 720
rect -624 708 -612 720
rect -600 708 -588 720
rect -576 708 -564 720
rect -552 708 -540 720
rect -528 708 -516 720
rect -504 708 -492 720
rect -480 708 -468 720
rect -456 708 -444 720
rect -432 708 -420 720
rect -408 708 -396 720
rect -384 708 -372 720
rect -360 708 -348 720
rect -336 708 -324 720
rect -312 708 -300 720
rect -288 708 -276 720
rect -264 708 -252 720
rect -240 708 -228 720
rect -216 708 -204 720
rect -192 708 -180 720
rect -168 708 -156 720
rect -144 708 -132 720
rect -120 708 -108 720
rect -96 708 -84 720
rect -72 708 -60 720
rect -48 708 -36 720
rect -24 708 -12 720
rect 0 708 12 720
rect 24 708 36 720
rect 48 708 60 720
rect 72 708 84 720
rect 96 708 108 720
rect 120 708 132 720
rect 144 708 156 720
rect 168 708 180 720
rect 192 708 204 720
rect 216 708 228 720
rect 240 708 252 720
rect 264 708 276 720
rect 288 708 300 720
rect 312 708 324 720
rect 336 708 348 720
rect 360 708 372 720
rect 384 708 396 720
rect 408 708 420 720
rect 432 708 444 720
rect 456 708 468 720
rect 480 708 492 720
rect 504 708 516 720
rect 528 708 540 720
rect 552 708 564 720
rect 576 708 588 720
rect 600 708 612 720
rect 624 708 636 720
rect 648 708 660 720
rect 672 708 684 720
rect 696 708 708 720
rect 720 708 732 720
rect 744 708 756 720
rect 768 708 780 720
rect 792 708 804 720
rect 816 708 828 720
rect 840 708 852 720
rect 864 708 876 720
rect 888 708 900 720
rect 912 708 924 720
rect 936 708 948 720
rect 960 708 972 720
rect 984 708 996 720
rect 1008 708 1020 720
rect 1032 708 1044 720
rect 1056 708 1068 720
rect 1080 708 1092 720
rect 1104 708 1116 720
rect 1128 708 1140 720
rect 1152 708 1164 720
rect 1176 708 1188 720
rect 1200 708 1212 720
rect 1224 708 1236 720
rect 1248 708 1260 720
rect 1272 708 1284 720
rect 1296 708 1308 720
rect 1320 708 1332 720
rect 1344 708 1356 720
rect 1368 708 1380 720
rect 1392 708 1404 720
rect 1416 708 1428 720
rect 1440 708 1452 720
rect 1464 708 1476 720
rect 1488 708 1500 720
rect 1512 708 1524 720
rect 1536 708 1548 720
rect 1560 708 1572 720
rect 1584 708 1596 720
rect 1608 708 1620 720
rect 1632 708 1644 720
rect 1656 708 1668 720
rect 1680 708 1692 720
rect 1704 708 1716 720
rect 1728 708 1740 720
rect 1752 708 1764 720
rect 1776 708 1788 720
rect 1800 708 1812 720
rect 1824 708 1836 720
rect 1848 708 1860 720
rect 1872 708 1884 720
rect 1896 708 1908 720
rect 1920 708 1932 720
rect 1944 708 1956 720
rect 1968 708 1980 720
rect 1992 708 2004 720
rect 2016 708 2028 720
rect 2040 708 2052 720
rect 2064 708 2076 720
rect 2088 708 2100 720
rect 2112 708 2124 720
rect 2136 708 2148 720
rect 2160 708 2172 720
rect 2184 708 2196 720
rect 2208 708 2220 720
rect 2232 708 2244 720
rect 2256 708 2268 720
rect 2280 708 2292 720
rect 2304 708 2316 720
rect 2328 708 2340 720
rect 2352 708 2364 720
rect 2376 708 2388 720
rect 2400 708 2412 720
rect 2424 708 2436 720
rect 2448 708 2460 720
rect 2472 708 2484 720
rect 2496 708 2508 720
rect 2520 708 2532 720
rect 2544 708 2556 720
rect 2568 708 2580 720
rect 2592 708 2604 720
rect 2616 708 2628 720
rect 2640 708 2652 720
rect 2664 708 2676 720
rect 2688 708 2700 720
rect 2712 708 2724 720
rect 2736 708 2748 720
rect 2760 708 2772 720
rect 2784 708 2796 720
rect 2808 708 2820 720
rect 2832 708 2844 720
rect 2856 708 2868 720
rect 2880 708 2892 720
rect 2904 708 2916 720
rect 2928 708 2940 720
rect 2952 708 2976 720
rect -1008 684 2976 708
rect -1008 672 -996 684
rect -984 672 -972 684
rect -960 672 -948 684
rect -936 672 -924 684
rect -912 672 -900 684
rect -888 672 -876 684
rect -864 672 -852 684
rect -840 672 -828 684
rect -816 672 -804 684
rect -792 672 -780 684
rect -768 672 -756 684
rect -744 672 -732 684
rect -720 672 -708 684
rect -696 672 -684 684
rect -672 672 -660 684
rect -648 672 -636 684
rect -624 672 -612 684
rect -600 672 -588 684
rect -576 672 -564 684
rect -552 672 -540 684
rect -528 672 -516 684
rect -504 672 -492 684
rect -480 672 -468 684
rect -456 672 -444 684
rect -432 672 -420 684
rect -408 672 -396 684
rect -384 672 -372 684
rect -360 672 -348 684
rect -336 672 -324 684
rect -312 672 -300 684
rect -288 672 -276 684
rect -264 672 -252 684
rect -240 672 -228 684
rect -216 672 -204 684
rect -192 672 -180 684
rect -168 672 -156 684
rect -144 672 -132 684
rect -120 672 -108 684
rect -96 672 -84 684
rect -72 672 -60 684
rect -48 672 -36 684
rect -24 672 -12 684
rect 0 672 12 684
rect 24 672 36 684
rect 48 672 60 684
rect 72 672 84 684
rect 96 672 108 684
rect 120 672 132 684
rect 144 672 156 684
rect 168 672 180 684
rect 192 672 204 684
rect 216 672 228 684
rect 240 672 252 684
rect 264 672 276 684
rect 288 672 300 684
rect 312 672 324 684
rect 336 672 348 684
rect 360 672 372 684
rect 384 672 396 684
rect 408 672 420 684
rect 432 672 444 684
rect 456 672 468 684
rect 480 672 492 684
rect 504 672 516 684
rect 528 672 540 684
rect 552 672 564 684
rect 576 672 588 684
rect 600 672 612 684
rect 624 672 636 684
rect 648 672 660 684
rect 672 672 684 684
rect 696 672 708 684
rect 720 672 732 684
rect 744 672 756 684
rect 768 672 780 684
rect 792 672 804 684
rect 816 672 828 684
rect 840 672 852 684
rect 864 672 876 684
rect 888 672 900 684
rect 912 672 924 684
rect 936 672 948 684
rect 960 672 972 684
rect 984 672 996 684
rect 1008 672 1020 684
rect 1032 672 1044 684
rect 1056 672 1068 684
rect 1080 672 1092 684
rect 1104 672 1116 684
rect 1128 672 1140 684
rect 1152 672 1164 684
rect 1176 672 1188 684
rect 1200 672 1212 684
rect 1224 672 1236 684
rect 1248 672 1260 684
rect 1272 672 1284 684
rect 1296 672 1308 684
rect 1320 672 1332 684
rect 1344 672 1356 684
rect 1368 672 1380 684
rect 1392 672 1404 684
rect 1416 672 1428 684
rect 1440 672 1452 684
rect 1464 672 1476 684
rect 1488 672 1500 684
rect 1512 672 1524 684
rect 1536 672 1548 684
rect 1560 672 1572 684
rect 1584 672 1596 684
rect 1608 672 1620 684
rect 1632 672 1644 684
rect 1656 672 1668 684
rect 1680 672 1692 684
rect 1704 672 1716 684
rect 1728 672 1740 684
rect 1752 672 1764 684
rect 1776 672 1788 684
rect 1800 672 1812 684
rect 1824 672 1836 684
rect 1848 672 1860 684
rect 1872 672 1884 684
rect 1896 672 1908 684
rect 1920 672 1932 684
rect 1944 672 1956 684
rect 1968 672 1980 684
rect 1992 672 2004 684
rect 2016 672 2028 684
rect 2040 672 2052 684
rect 2064 672 2076 684
rect 2088 672 2100 684
rect 2112 672 2124 684
rect 2136 672 2148 684
rect 2160 672 2172 684
rect 2184 672 2196 684
rect 2208 672 2220 684
rect 2232 672 2244 684
rect 2256 672 2268 684
rect 2280 672 2292 684
rect 2304 672 2316 684
rect 2328 672 2340 684
rect 2352 672 2364 684
rect 2376 672 2388 684
rect 2400 672 2412 684
rect 2424 672 2436 684
rect 2448 672 2460 684
rect 2472 672 2484 684
rect 2496 672 2508 684
rect 2520 672 2532 684
rect 2544 672 2556 684
rect 2568 672 2580 684
rect 2592 672 2604 684
rect 2616 672 2628 684
rect 2640 672 2652 684
rect 2664 672 2676 684
rect 2688 672 2700 684
rect 2712 672 2724 684
rect 2736 672 2748 684
rect 2760 672 2772 684
rect 2784 672 2796 684
rect 2808 672 2820 684
rect 2832 672 2844 684
rect 2856 672 2868 684
rect 2880 672 2892 684
rect 2904 672 2916 684
rect 2928 672 2940 684
rect 2952 672 2976 684
rect -1008 660 2976 672
rect -1008 -252 2976 -240
rect -1008 -264 -996 -252
rect -984 -264 -972 -252
rect -960 -264 -948 -252
rect -936 -264 -924 -252
rect -912 -264 -900 -252
rect -888 -264 -876 -252
rect -864 -264 -852 -252
rect -840 -264 -828 -252
rect -816 -264 -804 -252
rect -792 -264 -780 -252
rect -768 -264 -756 -252
rect -744 -264 -732 -252
rect -720 -264 -708 -252
rect -696 -264 -684 -252
rect -672 -264 -660 -252
rect -648 -264 -636 -252
rect -624 -264 -612 -252
rect -600 -264 -588 -252
rect -576 -264 -564 -252
rect -552 -264 -540 -252
rect -528 -264 -516 -252
rect -504 -264 -492 -252
rect -480 -264 -468 -252
rect -456 -264 -444 -252
rect -432 -264 -420 -252
rect -408 -264 -396 -252
rect -384 -264 -372 -252
rect -360 -264 -348 -252
rect -336 -264 -324 -252
rect -312 -264 -300 -252
rect -288 -264 -276 -252
rect -264 -264 -252 -252
rect -240 -264 -228 -252
rect -216 -264 -204 -252
rect -192 -264 -180 -252
rect -168 -264 -156 -252
rect -144 -264 -132 -252
rect -120 -264 -108 -252
rect -96 -264 -84 -252
rect -72 -264 -60 -252
rect -48 -264 -36 -252
rect -24 -264 -12 -252
rect 0 -264 12 -252
rect 24 -264 36 -252
rect 48 -264 60 -252
rect 72 -264 84 -252
rect 96 -264 108 -252
rect 120 -264 132 -252
rect 144 -264 156 -252
rect 168 -264 180 -252
rect 192 -264 204 -252
rect 216 -264 228 -252
rect 240 -264 252 -252
rect 264 -264 276 -252
rect 288 -264 300 -252
rect 312 -264 324 -252
rect 336 -264 348 -252
rect 360 -264 372 -252
rect 384 -264 396 -252
rect 408 -264 420 -252
rect 432 -264 444 -252
rect 456 -264 468 -252
rect 480 -264 492 -252
rect 504 -264 516 -252
rect 528 -264 540 -252
rect 552 -264 564 -252
rect 576 -264 588 -252
rect 600 -264 612 -252
rect 624 -264 636 -252
rect 648 -264 660 -252
rect 672 -264 684 -252
rect 696 -264 708 -252
rect 720 -264 732 -252
rect 744 -264 756 -252
rect 768 -264 780 -252
rect 792 -264 804 -252
rect 816 -264 828 -252
rect 840 -264 852 -252
rect 864 -264 876 -252
rect 888 -264 900 -252
rect 912 -264 924 -252
rect 936 -264 948 -252
rect 960 -264 972 -252
rect 984 -264 996 -252
rect 1008 -264 1020 -252
rect 1032 -264 1044 -252
rect 1056 -264 1068 -252
rect 1080 -264 1092 -252
rect 1104 -264 1116 -252
rect 1128 -264 1140 -252
rect 1152 -264 1164 -252
rect 1176 -264 1188 -252
rect 1200 -264 1212 -252
rect 1224 -264 1236 -252
rect 1248 -264 1260 -252
rect 1272 -264 1284 -252
rect 1296 -264 1308 -252
rect 1320 -264 1332 -252
rect 1344 -264 1356 -252
rect 1368 -264 1380 -252
rect 1392 -264 1404 -252
rect 1416 -264 1428 -252
rect 1440 -264 1452 -252
rect 1464 -264 1476 -252
rect 1488 -264 1500 -252
rect 1512 -264 1524 -252
rect 1536 -264 1548 -252
rect 1560 -264 1572 -252
rect 1584 -264 1596 -252
rect 1608 -264 1620 -252
rect 1632 -264 1644 -252
rect 1656 -264 1668 -252
rect 1680 -264 1692 -252
rect 1704 -264 1716 -252
rect 1728 -264 1740 -252
rect 1752 -264 1764 -252
rect 1776 -264 1788 -252
rect 1800 -264 1812 -252
rect 1824 -264 1836 -252
rect 1848 -264 1860 -252
rect 1872 -264 1884 -252
rect 1896 -264 1908 -252
rect 1920 -264 1932 -252
rect 1944 -264 1956 -252
rect 1968 -264 1980 -252
rect 1992 -264 2004 -252
rect 2016 -264 2028 -252
rect 2040 -264 2052 -252
rect 2064 -264 2076 -252
rect 2088 -264 2100 -252
rect 2112 -264 2124 -252
rect 2136 -264 2148 -252
rect 2160 -264 2172 -252
rect 2184 -264 2196 -252
rect 2208 -264 2220 -252
rect 2232 -264 2244 -252
rect 2256 -264 2268 -252
rect 2280 -264 2292 -252
rect 2304 -264 2316 -252
rect 2328 -264 2340 -252
rect 2352 -264 2364 -252
rect 2376 -264 2388 -252
rect 2400 -264 2412 -252
rect 2424 -264 2436 -252
rect 2448 -264 2460 -252
rect 2472 -264 2484 -252
rect 2496 -264 2508 -252
rect 2520 -264 2532 -252
rect 2544 -264 2556 -252
rect 2568 -264 2580 -252
rect 2592 -264 2604 -252
rect 2616 -264 2628 -252
rect 2640 -264 2652 -252
rect 2664 -264 2676 -252
rect 2688 -264 2700 -252
rect 2712 -264 2724 -252
rect 2736 -264 2748 -252
rect 2760 -264 2772 -252
rect 2784 -264 2796 -252
rect 2808 -264 2820 -252
rect 2832 -264 2844 -252
rect 2856 -264 2868 -252
rect 2880 -264 2892 -252
rect 2904 -264 2916 -252
rect 2928 -264 2940 -252
rect 2952 -264 2976 -252
rect -1008 -288 2976 -264
rect -1008 -300 -996 -288
rect -984 -300 -972 -288
rect -960 -300 -948 -288
rect -936 -300 -924 -288
rect -912 -300 -900 -288
rect -888 -300 -876 -288
rect -864 -300 -852 -288
rect -840 -300 -828 -288
rect -816 -300 -804 -288
rect -792 -300 -780 -288
rect -768 -300 -756 -288
rect -744 -300 -732 -288
rect -720 -300 -708 -288
rect -696 -300 -684 -288
rect -672 -300 -660 -288
rect -648 -300 -636 -288
rect -624 -300 -612 -288
rect -600 -300 -588 -288
rect -576 -300 -564 -288
rect -552 -300 -540 -288
rect -528 -300 -516 -288
rect -504 -300 -492 -288
rect -480 -300 -468 -288
rect -456 -300 -444 -288
rect -432 -300 -420 -288
rect -408 -300 -396 -288
rect -384 -300 -372 -288
rect -360 -300 -348 -288
rect -336 -300 -324 -288
rect -312 -300 -300 -288
rect -288 -300 -276 -288
rect -264 -300 -252 -288
rect -240 -300 -228 -288
rect -216 -300 -204 -288
rect -192 -300 -180 -288
rect -168 -300 -156 -288
rect -144 -300 -132 -288
rect -120 -300 -108 -288
rect -96 -300 -84 -288
rect -72 -300 -60 -288
rect -48 -300 -36 -288
rect -24 -300 -12 -288
rect 0 -300 12 -288
rect 24 -300 36 -288
rect 48 -300 60 -288
rect 72 -300 84 -288
rect 96 -300 108 -288
rect 120 -300 132 -288
rect 144 -300 156 -288
rect 168 -300 180 -288
rect 192 -300 204 -288
rect 216 -300 228 -288
rect 240 -300 252 -288
rect 264 -300 276 -288
rect 288 -300 300 -288
rect 312 -300 324 -288
rect 336 -300 348 -288
rect 360 -300 372 -288
rect 384 -300 396 -288
rect 408 -300 420 -288
rect 432 -300 444 -288
rect 456 -300 468 -288
rect 480 -300 492 -288
rect 504 -300 516 -288
rect 528 -300 540 -288
rect 552 -300 564 -288
rect 576 -300 588 -288
rect 600 -300 612 -288
rect 624 -300 636 -288
rect 648 -300 660 -288
rect 672 -300 684 -288
rect 696 -300 708 -288
rect 720 -300 732 -288
rect 744 -300 756 -288
rect 768 -300 780 -288
rect 792 -300 804 -288
rect 816 -300 828 -288
rect 840 -300 852 -288
rect 864 -300 876 -288
rect 888 -300 900 -288
rect 912 -300 924 -288
rect 936 -300 948 -288
rect 960 -300 972 -288
rect 984 -300 996 -288
rect 1008 -300 1020 -288
rect 1032 -300 1044 -288
rect 1056 -300 1068 -288
rect 1080 -300 1092 -288
rect 1104 -300 1116 -288
rect 1128 -300 1140 -288
rect 1152 -300 1164 -288
rect 1176 -300 1188 -288
rect 1200 -300 1212 -288
rect 1224 -300 1236 -288
rect 1248 -300 1260 -288
rect 1272 -300 1284 -288
rect 1296 -300 1308 -288
rect 1320 -300 1332 -288
rect 1344 -300 1356 -288
rect 1368 -300 1380 -288
rect 1392 -300 1404 -288
rect 1416 -300 1428 -288
rect 1440 -300 1452 -288
rect 1464 -300 1476 -288
rect 1488 -300 1500 -288
rect 1512 -300 1524 -288
rect 1536 -300 1548 -288
rect 1560 -300 1572 -288
rect 1584 -300 1596 -288
rect 1608 -300 1620 -288
rect 1632 -300 1644 -288
rect 1656 -300 1668 -288
rect 1680 -300 1692 -288
rect 1704 -300 1716 -288
rect 1728 -300 1740 -288
rect 1752 -300 1764 -288
rect 1776 -300 1788 -288
rect 1800 -300 1812 -288
rect 1824 -300 1836 -288
rect 1848 -300 1860 -288
rect 1872 -300 1884 -288
rect 1896 -300 1908 -288
rect 1920 -300 1932 -288
rect 1944 -300 1956 -288
rect 1968 -300 1980 -288
rect 1992 -300 2004 -288
rect 2016 -300 2028 -288
rect 2040 -300 2052 -288
rect 2064 -300 2076 -288
rect 2088 -300 2100 -288
rect 2112 -300 2124 -288
rect 2136 -300 2148 -288
rect 2160 -300 2172 -288
rect 2184 -300 2196 -288
rect 2208 -300 2220 -288
rect 2232 -300 2244 -288
rect 2256 -300 2268 -288
rect 2280 -300 2292 -288
rect 2304 -300 2316 -288
rect 2328 -300 2340 -288
rect 2352 -300 2364 -288
rect 2376 -300 2388 -288
rect 2400 -300 2412 -288
rect 2424 -300 2436 -288
rect 2448 -300 2460 -288
rect 2472 -300 2484 -288
rect 2496 -300 2508 -288
rect 2520 -300 2532 -288
rect 2544 -300 2556 -288
rect 2568 -300 2580 -288
rect 2592 -300 2604 -288
rect 2616 -300 2628 -288
rect 2640 -300 2652 -288
rect 2664 -300 2676 -288
rect 2688 -300 2700 -288
rect 2712 -300 2724 -288
rect 2736 -300 2748 -288
rect 2760 -300 2772 -288
rect 2784 -300 2796 -288
rect 2808 -300 2820 -288
rect 2832 -300 2844 -288
rect 2856 -300 2868 -288
rect 2880 -300 2892 -288
rect 2904 -300 2916 -288
rect 2928 -300 2940 -288
rect 2952 -300 2976 -288
rect -1008 -324 2976 -300
rect -1008 -336 -996 -324
rect -984 -336 -972 -324
rect -960 -336 -948 -324
rect -936 -336 -924 -324
rect -912 -336 -900 -324
rect -888 -336 -876 -324
rect -864 -336 -852 -324
rect -840 -336 -828 -324
rect -816 -336 -804 -324
rect -792 -336 -780 -324
rect -768 -336 -756 -324
rect -744 -336 -732 -324
rect -720 -336 -708 -324
rect -696 -336 -684 -324
rect -672 -336 -660 -324
rect -648 -336 -636 -324
rect -624 -336 -612 -324
rect -600 -336 -588 -324
rect -576 -336 -564 -324
rect -552 -336 -540 -324
rect -528 -336 -516 -324
rect -504 -336 -492 -324
rect -480 -336 -468 -324
rect -456 -336 -444 -324
rect -432 -336 -420 -324
rect -408 -336 -396 -324
rect -384 -336 -372 -324
rect -360 -336 -348 -324
rect -336 -336 -324 -324
rect -312 -336 -300 -324
rect -288 -336 -276 -324
rect -264 -336 -252 -324
rect -240 -336 -228 -324
rect -216 -336 -204 -324
rect -192 -336 -180 -324
rect -168 -336 -156 -324
rect -144 -336 -132 -324
rect -120 -336 -108 -324
rect -96 -336 -84 -324
rect -72 -336 -60 -324
rect -48 -336 -36 -324
rect -24 -336 -12 -324
rect 0 -336 12 -324
rect 24 -336 36 -324
rect 48 -336 60 -324
rect 72 -336 84 -324
rect 96 -336 108 -324
rect 120 -336 132 -324
rect 144 -336 156 -324
rect 168 -336 180 -324
rect 192 -336 204 -324
rect 216 -336 228 -324
rect 240 -336 252 -324
rect 264 -336 276 -324
rect 288 -336 300 -324
rect 312 -336 324 -324
rect 336 -336 348 -324
rect 360 -336 372 -324
rect 384 -336 396 -324
rect 408 -336 420 -324
rect 432 -336 444 -324
rect 456 -336 468 -324
rect 480 -336 492 -324
rect 504 -336 516 -324
rect 528 -336 540 -324
rect 552 -336 564 -324
rect 576 -336 588 -324
rect 600 -336 612 -324
rect 624 -336 636 -324
rect 648 -336 660 -324
rect 672 -336 684 -324
rect 696 -336 708 -324
rect 720 -336 732 -324
rect 744 -336 756 -324
rect 768 -336 780 -324
rect 792 -336 804 -324
rect 816 -336 828 -324
rect 840 -336 852 -324
rect 864 -336 876 -324
rect 888 -336 900 -324
rect 912 -336 924 -324
rect 936 -336 948 -324
rect 960 -336 972 -324
rect 984 -336 996 -324
rect 1008 -336 1020 -324
rect 1032 -336 1044 -324
rect 1056 -336 1068 -324
rect 1080 -336 1092 -324
rect 1104 -336 1116 -324
rect 1128 -336 1140 -324
rect 1152 -336 1164 -324
rect 1176 -336 1188 -324
rect 1200 -336 1212 -324
rect 1224 -336 1236 -324
rect 1248 -336 1260 -324
rect 1272 -336 1284 -324
rect 1296 -336 1308 -324
rect 1320 -336 1332 -324
rect 1344 -336 1356 -324
rect 1368 -336 1380 -324
rect 1392 -336 1404 -324
rect 1416 -336 1428 -324
rect 1440 -336 1452 -324
rect 1464 -336 1476 -324
rect 1488 -336 1500 -324
rect 1512 -336 1524 -324
rect 1536 -336 1548 -324
rect 1560 -336 1572 -324
rect 1584 -336 1596 -324
rect 1608 -336 1620 -324
rect 1632 -336 1644 -324
rect 1656 -336 1668 -324
rect 1680 -336 1692 -324
rect 1704 -336 1716 -324
rect 1728 -336 1740 -324
rect 1752 -336 1764 -324
rect 1776 -336 1788 -324
rect 1800 -336 1812 -324
rect 1824 -336 1836 -324
rect 1848 -336 1860 -324
rect 1872 -336 1884 -324
rect 1896 -336 1908 -324
rect 1920 -336 1932 -324
rect 1944 -336 1956 -324
rect 1968 -336 1980 -324
rect 1992 -336 2004 -324
rect 2016 -336 2028 -324
rect 2040 -336 2052 -324
rect 2064 -336 2076 -324
rect 2088 -336 2100 -324
rect 2112 -336 2124 -324
rect 2136 -336 2148 -324
rect 2160 -336 2172 -324
rect 2184 -336 2196 -324
rect 2208 -336 2220 -324
rect 2232 -336 2244 -324
rect 2256 -336 2268 -324
rect 2280 -336 2292 -324
rect 2304 -336 2316 -324
rect 2328 -336 2340 -324
rect 2352 -336 2364 -324
rect 2376 -336 2388 -324
rect 2400 -336 2412 -324
rect 2424 -336 2436 -324
rect 2448 -336 2460 -324
rect 2472 -336 2484 -324
rect 2496 -336 2508 -324
rect 2520 -336 2532 -324
rect 2544 -336 2556 -324
rect 2568 -336 2580 -324
rect 2592 -336 2604 -324
rect 2616 -336 2628 -324
rect 2640 -336 2652 -324
rect 2664 -336 2676 -324
rect 2688 -336 2700 -324
rect 2712 -336 2724 -324
rect 2736 -336 2748 -324
rect 2760 -336 2772 -324
rect 2784 -336 2796 -324
rect 2808 -336 2820 -324
rect 2832 -336 2844 -324
rect 2856 -336 2868 -324
rect 2880 -336 2892 -324
rect 2904 -336 2916 -324
rect 2928 -336 2940 -324
rect 2952 -336 2976 -324
rect -1008 -360 2976 -336
rect -1008 -372 -996 -360
rect -984 -372 -972 -360
rect -960 -372 -948 -360
rect -936 -372 -924 -360
rect -912 -372 -900 -360
rect -888 -372 -876 -360
rect -864 -372 -852 -360
rect -840 -372 -828 -360
rect -816 -372 -804 -360
rect -792 -372 -780 -360
rect -768 -372 -756 -360
rect -744 -372 -732 -360
rect -720 -372 -708 -360
rect -696 -372 -684 -360
rect -672 -372 -660 -360
rect -648 -372 -636 -360
rect -624 -372 -612 -360
rect -600 -372 -588 -360
rect -576 -372 -564 -360
rect -552 -372 -540 -360
rect -528 -372 -516 -360
rect -504 -372 -492 -360
rect -480 -372 -468 -360
rect -456 -372 -444 -360
rect -432 -372 -420 -360
rect -408 -372 -396 -360
rect -384 -372 -372 -360
rect -360 -372 -348 -360
rect -336 -372 -324 -360
rect -312 -372 -300 -360
rect -288 -372 -276 -360
rect -264 -372 -252 -360
rect -240 -372 -228 -360
rect -216 -372 -204 -360
rect -192 -372 -180 -360
rect -168 -372 -156 -360
rect -144 -372 -132 -360
rect -120 -372 -108 -360
rect -96 -372 -84 -360
rect -72 -372 -60 -360
rect -48 -372 -36 -360
rect -24 -372 -12 -360
rect 0 -372 12 -360
rect 24 -372 36 -360
rect 48 -372 60 -360
rect 72 -372 84 -360
rect 96 -372 108 -360
rect 120 -372 132 -360
rect 144 -372 156 -360
rect 168 -372 180 -360
rect 192 -372 204 -360
rect 216 -372 228 -360
rect 240 -372 252 -360
rect 264 -372 276 -360
rect 288 -372 300 -360
rect 312 -372 324 -360
rect 336 -372 348 -360
rect 360 -372 372 -360
rect 384 -372 396 -360
rect 408 -372 420 -360
rect 432 -372 444 -360
rect 456 -372 468 -360
rect 480 -372 492 -360
rect 504 -372 516 -360
rect 528 -372 540 -360
rect 552 -372 564 -360
rect 576 -372 588 -360
rect 600 -372 612 -360
rect 624 -372 636 -360
rect 648 -372 660 -360
rect 672 -372 684 -360
rect 696 -372 708 -360
rect 720 -372 732 -360
rect 744 -372 756 -360
rect 768 -372 780 -360
rect 792 -372 804 -360
rect 816 -372 828 -360
rect 840 -372 852 -360
rect 864 -372 876 -360
rect 888 -372 900 -360
rect 912 -372 924 -360
rect 936 -372 948 -360
rect 960 -372 972 -360
rect 984 -372 996 -360
rect 1008 -372 1020 -360
rect 1032 -372 1044 -360
rect 1056 -372 1068 -360
rect 1080 -372 1092 -360
rect 1104 -372 1116 -360
rect 1128 -372 1140 -360
rect 1152 -372 1164 -360
rect 1176 -372 1188 -360
rect 1200 -372 1212 -360
rect 1224 -372 1236 -360
rect 1248 -372 1260 -360
rect 1272 -372 1284 -360
rect 1296 -372 1308 -360
rect 1320 -372 1332 -360
rect 1344 -372 1356 -360
rect 1368 -372 1380 -360
rect 1392 -372 1404 -360
rect 1416 -372 1428 -360
rect 1440 -372 1452 -360
rect 1464 -372 1476 -360
rect 1488 -372 1500 -360
rect 1512 -372 1524 -360
rect 1536 -372 1548 -360
rect 1560 -372 1572 -360
rect 1584 -372 1596 -360
rect 1608 -372 1620 -360
rect 1632 -372 1644 -360
rect 1656 -372 1668 -360
rect 1680 -372 1692 -360
rect 1704 -372 1716 -360
rect 1728 -372 1740 -360
rect 1752 -372 1764 -360
rect 1776 -372 1788 -360
rect 1800 -372 1812 -360
rect 1824 -372 1836 -360
rect 1848 -372 1860 -360
rect 1872 -372 1884 -360
rect 1896 -372 1908 -360
rect 1920 -372 1932 -360
rect 1944 -372 1956 -360
rect 1968 -372 1980 -360
rect 1992 -372 2004 -360
rect 2016 -372 2028 -360
rect 2040 -372 2052 -360
rect 2064 -372 2076 -360
rect 2088 -372 2100 -360
rect 2112 -372 2124 -360
rect 2136 -372 2148 -360
rect 2160 -372 2172 -360
rect 2184 -372 2196 -360
rect 2208 -372 2220 -360
rect 2232 -372 2244 -360
rect 2256 -372 2268 -360
rect 2280 -372 2292 -360
rect 2304 -372 2316 -360
rect 2328 -372 2340 -360
rect 2352 -372 2364 -360
rect 2376 -372 2388 -360
rect 2400 -372 2412 -360
rect 2424 -372 2436 -360
rect 2448 -372 2460 -360
rect 2472 -372 2484 -360
rect 2496 -372 2508 -360
rect 2520 -372 2532 -360
rect 2544 -372 2556 -360
rect 2568 -372 2580 -360
rect 2592 -372 2604 -360
rect 2616 -372 2628 -360
rect 2640 -372 2652 -360
rect 2664 -372 2676 -360
rect 2688 -372 2700 -360
rect 2712 -372 2724 -360
rect 2736 -372 2748 -360
rect 2760 -372 2772 -360
rect 2784 -372 2796 -360
rect 2808 -372 2820 -360
rect 2832 -372 2844 -360
rect 2856 -372 2868 -360
rect 2880 -372 2892 -360
rect 2904 -372 2916 -360
rect 2928 -372 2940 -360
rect 2952 -372 2976 -360
rect -1008 -384 2976 -372
<< mimcapcontact >>
rect -996 780 -984 792
rect -972 780 -960 792
rect -948 780 -936 792
rect -924 780 -912 792
rect -900 780 -888 792
rect -876 780 -864 792
rect -852 780 -840 792
rect -828 780 -816 792
rect -804 780 -792 792
rect -780 780 -768 792
rect -756 780 -744 792
rect -732 780 -720 792
rect -708 780 -696 792
rect -684 780 -672 792
rect -660 780 -648 792
rect -636 780 -624 792
rect -612 780 -600 792
rect -588 780 -576 792
rect -564 780 -552 792
rect -540 780 -528 792
rect -516 780 -504 792
rect -492 780 -480 792
rect -468 780 -456 792
rect -444 780 -432 792
rect -420 780 -408 792
rect -396 780 -384 792
rect -372 780 -360 792
rect -348 780 -336 792
rect -324 780 -312 792
rect -300 780 -288 792
rect -276 780 -264 792
rect -252 780 -240 792
rect -228 780 -216 792
rect -204 780 -192 792
rect -180 780 -168 792
rect -156 780 -144 792
rect -132 780 -120 792
rect -108 780 -96 792
rect -84 780 -72 792
rect -60 780 -48 792
rect -36 780 -24 792
rect -12 780 0 792
rect 12 780 24 792
rect 36 780 48 792
rect 60 780 72 792
rect 84 780 96 792
rect 108 780 120 792
rect 132 780 144 792
rect 156 780 168 792
rect 180 780 192 792
rect 204 780 216 792
rect 228 780 240 792
rect 252 780 264 792
rect 276 780 288 792
rect 300 780 312 792
rect 324 780 336 792
rect 348 780 360 792
rect 372 780 384 792
rect 396 780 408 792
rect 420 780 432 792
rect 444 780 456 792
rect 468 780 480 792
rect 492 780 504 792
rect 516 780 528 792
rect 540 780 552 792
rect 564 780 576 792
rect 588 780 600 792
rect 612 780 624 792
rect 636 780 648 792
rect 660 780 672 792
rect 684 780 696 792
rect 708 780 720 792
rect 732 780 744 792
rect 756 780 768 792
rect 780 780 792 792
rect 804 780 816 792
rect 828 780 840 792
rect 852 780 864 792
rect 876 780 888 792
rect 900 780 912 792
rect 924 780 936 792
rect 948 780 960 792
rect 972 780 984 792
rect 996 780 1008 792
rect 1020 780 1032 792
rect 1044 780 1056 792
rect 1068 780 1080 792
rect 1092 780 1104 792
rect 1116 780 1128 792
rect 1140 780 1152 792
rect 1164 780 1176 792
rect 1188 780 1200 792
rect 1212 780 1224 792
rect 1236 780 1248 792
rect 1260 780 1272 792
rect 1284 780 1296 792
rect 1308 780 1320 792
rect 1332 780 1344 792
rect 1356 780 1368 792
rect 1380 780 1392 792
rect 1404 780 1416 792
rect 1428 780 1440 792
rect 1452 780 1464 792
rect 1476 780 1488 792
rect 1500 780 1512 792
rect 1524 780 1536 792
rect 1548 780 1560 792
rect 1572 780 1584 792
rect 1596 780 1608 792
rect 1620 780 1632 792
rect 1644 780 1656 792
rect 1668 780 1680 792
rect 1692 780 1704 792
rect 1716 780 1728 792
rect 1740 780 1752 792
rect 1764 780 1776 792
rect 1788 780 1800 792
rect 1812 780 1824 792
rect 1836 780 1848 792
rect 1860 780 1872 792
rect 1884 780 1896 792
rect 1908 780 1920 792
rect 1932 780 1944 792
rect 1956 780 1968 792
rect 1980 780 1992 792
rect 2004 780 2016 792
rect 2028 780 2040 792
rect 2052 780 2064 792
rect 2076 780 2088 792
rect 2100 780 2112 792
rect 2124 780 2136 792
rect 2148 780 2160 792
rect 2172 780 2184 792
rect 2196 780 2208 792
rect 2220 780 2232 792
rect 2244 780 2256 792
rect 2268 780 2280 792
rect 2292 780 2304 792
rect 2316 780 2328 792
rect 2340 780 2352 792
rect 2364 780 2376 792
rect 2388 780 2400 792
rect 2412 780 2424 792
rect 2436 780 2448 792
rect 2460 780 2472 792
rect 2484 780 2496 792
rect 2508 780 2520 792
rect 2532 780 2544 792
rect 2556 780 2568 792
rect 2580 780 2592 792
rect 2604 780 2616 792
rect 2628 780 2640 792
rect 2652 780 2664 792
rect 2676 780 2688 792
rect 2700 780 2712 792
rect 2724 780 2736 792
rect 2748 780 2760 792
rect 2772 780 2784 792
rect 2796 780 2808 792
rect 2820 780 2832 792
rect 2844 780 2856 792
rect 2868 780 2880 792
rect 2892 780 2904 792
rect 2916 780 2928 792
rect 2940 780 2952 792
rect -996 744 -984 756
rect -972 744 -960 756
rect -948 744 -936 756
rect -924 744 -912 756
rect -900 744 -888 756
rect -876 744 -864 756
rect -852 744 -840 756
rect -828 744 -816 756
rect -804 744 -792 756
rect -780 744 -768 756
rect -756 744 -744 756
rect -732 744 -720 756
rect -708 744 -696 756
rect -684 744 -672 756
rect -660 744 -648 756
rect -636 744 -624 756
rect -612 744 -600 756
rect -588 744 -576 756
rect -564 744 -552 756
rect -540 744 -528 756
rect -516 744 -504 756
rect -492 744 -480 756
rect -468 744 -456 756
rect -444 744 -432 756
rect -420 744 -408 756
rect -396 744 -384 756
rect -372 744 -360 756
rect -348 744 -336 756
rect -324 744 -312 756
rect -300 744 -288 756
rect -276 744 -264 756
rect -252 744 -240 756
rect -228 744 -216 756
rect -204 744 -192 756
rect -180 744 -168 756
rect -156 744 -144 756
rect -132 744 -120 756
rect -108 744 -96 756
rect -84 744 -72 756
rect -60 744 -48 756
rect -36 744 -24 756
rect -12 744 0 756
rect 12 744 24 756
rect 36 744 48 756
rect 60 744 72 756
rect 84 744 96 756
rect 108 744 120 756
rect 132 744 144 756
rect 156 744 168 756
rect 180 744 192 756
rect 204 744 216 756
rect 228 744 240 756
rect 252 744 264 756
rect 276 744 288 756
rect 300 744 312 756
rect 324 744 336 756
rect 348 744 360 756
rect 372 744 384 756
rect 396 744 408 756
rect 420 744 432 756
rect 444 744 456 756
rect 468 744 480 756
rect 492 744 504 756
rect 516 744 528 756
rect 540 744 552 756
rect 564 744 576 756
rect 588 744 600 756
rect 612 744 624 756
rect 636 744 648 756
rect 660 744 672 756
rect 684 744 696 756
rect 708 744 720 756
rect 732 744 744 756
rect 756 744 768 756
rect 780 744 792 756
rect 804 744 816 756
rect 828 744 840 756
rect 852 744 864 756
rect 876 744 888 756
rect 900 744 912 756
rect 924 744 936 756
rect 948 744 960 756
rect 972 744 984 756
rect 996 744 1008 756
rect 1020 744 1032 756
rect 1044 744 1056 756
rect 1068 744 1080 756
rect 1092 744 1104 756
rect 1116 744 1128 756
rect 1140 744 1152 756
rect 1164 744 1176 756
rect 1188 744 1200 756
rect 1212 744 1224 756
rect 1236 744 1248 756
rect 1260 744 1272 756
rect 1284 744 1296 756
rect 1308 744 1320 756
rect 1332 744 1344 756
rect 1356 744 1368 756
rect 1380 744 1392 756
rect 1404 744 1416 756
rect 1428 744 1440 756
rect 1452 744 1464 756
rect 1476 744 1488 756
rect 1500 744 1512 756
rect 1524 744 1536 756
rect 1548 744 1560 756
rect 1572 744 1584 756
rect 1596 744 1608 756
rect 1620 744 1632 756
rect 1644 744 1656 756
rect 1668 744 1680 756
rect 1692 744 1704 756
rect 1716 744 1728 756
rect 1740 744 1752 756
rect 1764 744 1776 756
rect 1788 744 1800 756
rect 1812 744 1824 756
rect 1836 744 1848 756
rect 1860 744 1872 756
rect 1884 744 1896 756
rect 1908 744 1920 756
rect 1932 744 1944 756
rect 1956 744 1968 756
rect 1980 744 1992 756
rect 2004 744 2016 756
rect 2028 744 2040 756
rect 2052 744 2064 756
rect 2076 744 2088 756
rect 2100 744 2112 756
rect 2124 744 2136 756
rect 2148 744 2160 756
rect 2172 744 2184 756
rect 2196 744 2208 756
rect 2220 744 2232 756
rect 2244 744 2256 756
rect 2268 744 2280 756
rect 2292 744 2304 756
rect 2316 744 2328 756
rect 2340 744 2352 756
rect 2364 744 2376 756
rect 2388 744 2400 756
rect 2412 744 2424 756
rect 2436 744 2448 756
rect 2460 744 2472 756
rect 2484 744 2496 756
rect 2508 744 2520 756
rect 2532 744 2544 756
rect 2556 744 2568 756
rect 2580 744 2592 756
rect 2604 744 2616 756
rect 2628 744 2640 756
rect 2652 744 2664 756
rect 2676 744 2688 756
rect 2700 744 2712 756
rect 2724 744 2736 756
rect 2748 744 2760 756
rect 2772 744 2784 756
rect 2796 744 2808 756
rect 2820 744 2832 756
rect 2844 744 2856 756
rect 2868 744 2880 756
rect 2892 744 2904 756
rect 2916 744 2928 756
rect 2940 744 2952 756
rect -996 708 -984 720
rect -972 708 -960 720
rect -948 708 -936 720
rect -924 708 -912 720
rect -900 708 -888 720
rect -876 708 -864 720
rect -852 708 -840 720
rect -828 708 -816 720
rect -804 708 -792 720
rect -780 708 -768 720
rect -756 708 -744 720
rect -732 708 -720 720
rect -708 708 -696 720
rect -684 708 -672 720
rect -660 708 -648 720
rect -636 708 -624 720
rect -612 708 -600 720
rect -588 708 -576 720
rect -564 708 -552 720
rect -540 708 -528 720
rect -516 708 -504 720
rect -492 708 -480 720
rect -468 708 -456 720
rect -444 708 -432 720
rect -420 708 -408 720
rect -396 708 -384 720
rect -372 708 -360 720
rect -348 708 -336 720
rect -324 708 -312 720
rect -300 708 -288 720
rect -276 708 -264 720
rect -252 708 -240 720
rect -228 708 -216 720
rect -204 708 -192 720
rect -180 708 -168 720
rect -156 708 -144 720
rect -132 708 -120 720
rect -108 708 -96 720
rect -84 708 -72 720
rect -60 708 -48 720
rect -36 708 -24 720
rect -12 708 0 720
rect 12 708 24 720
rect 36 708 48 720
rect 60 708 72 720
rect 84 708 96 720
rect 108 708 120 720
rect 132 708 144 720
rect 156 708 168 720
rect 180 708 192 720
rect 204 708 216 720
rect 228 708 240 720
rect 252 708 264 720
rect 276 708 288 720
rect 300 708 312 720
rect 324 708 336 720
rect 348 708 360 720
rect 372 708 384 720
rect 396 708 408 720
rect 420 708 432 720
rect 444 708 456 720
rect 468 708 480 720
rect 492 708 504 720
rect 516 708 528 720
rect 540 708 552 720
rect 564 708 576 720
rect 588 708 600 720
rect 612 708 624 720
rect 636 708 648 720
rect 660 708 672 720
rect 684 708 696 720
rect 708 708 720 720
rect 732 708 744 720
rect 756 708 768 720
rect 780 708 792 720
rect 804 708 816 720
rect 828 708 840 720
rect 852 708 864 720
rect 876 708 888 720
rect 900 708 912 720
rect 924 708 936 720
rect 948 708 960 720
rect 972 708 984 720
rect 996 708 1008 720
rect 1020 708 1032 720
rect 1044 708 1056 720
rect 1068 708 1080 720
rect 1092 708 1104 720
rect 1116 708 1128 720
rect 1140 708 1152 720
rect 1164 708 1176 720
rect 1188 708 1200 720
rect 1212 708 1224 720
rect 1236 708 1248 720
rect 1260 708 1272 720
rect 1284 708 1296 720
rect 1308 708 1320 720
rect 1332 708 1344 720
rect 1356 708 1368 720
rect 1380 708 1392 720
rect 1404 708 1416 720
rect 1428 708 1440 720
rect 1452 708 1464 720
rect 1476 708 1488 720
rect 1500 708 1512 720
rect 1524 708 1536 720
rect 1548 708 1560 720
rect 1572 708 1584 720
rect 1596 708 1608 720
rect 1620 708 1632 720
rect 1644 708 1656 720
rect 1668 708 1680 720
rect 1692 708 1704 720
rect 1716 708 1728 720
rect 1740 708 1752 720
rect 1764 708 1776 720
rect 1788 708 1800 720
rect 1812 708 1824 720
rect 1836 708 1848 720
rect 1860 708 1872 720
rect 1884 708 1896 720
rect 1908 708 1920 720
rect 1932 708 1944 720
rect 1956 708 1968 720
rect 1980 708 1992 720
rect 2004 708 2016 720
rect 2028 708 2040 720
rect 2052 708 2064 720
rect 2076 708 2088 720
rect 2100 708 2112 720
rect 2124 708 2136 720
rect 2148 708 2160 720
rect 2172 708 2184 720
rect 2196 708 2208 720
rect 2220 708 2232 720
rect 2244 708 2256 720
rect 2268 708 2280 720
rect 2292 708 2304 720
rect 2316 708 2328 720
rect 2340 708 2352 720
rect 2364 708 2376 720
rect 2388 708 2400 720
rect 2412 708 2424 720
rect 2436 708 2448 720
rect 2460 708 2472 720
rect 2484 708 2496 720
rect 2508 708 2520 720
rect 2532 708 2544 720
rect 2556 708 2568 720
rect 2580 708 2592 720
rect 2604 708 2616 720
rect 2628 708 2640 720
rect 2652 708 2664 720
rect 2676 708 2688 720
rect 2700 708 2712 720
rect 2724 708 2736 720
rect 2748 708 2760 720
rect 2772 708 2784 720
rect 2796 708 2808 720
rect 2820 708 2832 720
rect 2844 708 2856 720
rect 2868 708 2880 720
rect 2892 708 2904 720
rect 2916 708 2928 720
rect 2940 708 2952 720
rect -996 672 -984 684
rect -972 672 -960 684
rect -948 672 -936 684
rect -924 672 -912 684
rect -900 672 -888 684
rect -876 672 -864 684
rect -852 672 -840 684
rect -828 672 -816 684
rect -804 672 -792 684
rect -780 672 -768 684
rect -756 672 -744 684
rect -732 672 -720 684
rect -708 672 -696 684
rect -684 672 -672 684
rect -660 672 -648 684
rect -636 672 -624 684
rect -612 672 -600 684
rect -588 672 -576 684
rect -564 672 -552 684
rect -540 672 -528 684
rect -516 672 -504 684
rect -492 672 -480 684
rect -468 672 -456 684
rect -444 672 -432 684
rect -420 672 -408 684
rect -396 672 -384 684
rect -372 672 -360 684
rect -348 672 -336 684
rect -324 672 -312 684
rect -300 672 -288 684
rect -276 672 -264 684
rect -252 672 -240 684
rect -228 672 -216 684
rect -204 672 -192 684
rect -180 672 -168 684
rect -156 672 -144 684
rect -132 672 -120 684
rect -108 672 -96 684
rect -84 672 -72 684
rect -60 672 -48 684
rect -36 672 -24 684
rect -12 672 0 684
rect 12 672 24 684
rect 36 672 48 684
rect 60 672 72 684
rect 84 672 96 684
rect 108 672 120 684
rect 132 672 144 684
rect 156 672 168 684
rect 180 672 192 684
rect 204 672 216 684
rect 228 672 240 684
rect 252 672 264 684
rect 276 672 288 684
rect 300 672 312 684
rect 324 672 336 684
rect 348 672 360 684
rect 372 672 384 684
rect 396 672 408 684
rect 420 672 432 684
rect 444 672 456 684
rect 468 672 480 684
rect 492 672 504 684
rect 516 672 528 684
rect 540 672 552 684
rect 564 672 576 684
rect 588 672 600 684
rect 612 672 624 684
rect 636 672 648 684
rect 660 672 672 684
rect 684 672 696 684
rect 708 672 720 684
rect 732 672 744 684
rect 756 672 768 684
rect 780 672 792 684
rect 804 672 816 684
rect 828 672 840 684
rect 852 672 864 684
rect 876 672 888 684
rect 900 672 912 684
rect 924 672 936 684
rect 948 672 960 684
rect 972 672 984 684
rect 996 672 1008 684
rect 1020 672 1032 684
rect 1044 672 1056 684
rect 1068 672 1080 684
rect 1092 672 1104 684
rect 1116 672 1128 684
rect 1140 672 1152 684
rect 1164 672 1176 684
rect 1188 672 1200 684
rect 1212 672 1224 684
rect 1236 672 1248 684
rect 1260 672 1272 684
rect 1284 672 1296 684
rect 1308 672 1320 684
rect 1332 672 1344 684
rect 1356 672 1368 684
rect 1380 672 1392 684
rect 1404 672 1416 684
rect 1428 672 1440 684
rect 1452 672 1464 684
rect 1476 672 1488 684
rect 1500 672 1512 684
rect 1524 672 1536 684
rect 1548 672 1560 684
rect 1572 672 1584 684
rect 1596 672 1608 684
rect 1620 672 1632 684
rect 1644 672 1656 684
rect 1668 672 1680 684
rect 1692 672 1704 684
rect 1716 672 1728 684
rect 1740 672 1752 684
rect 1764 672 1776 684
rect 1788 672 1800 684
rect 1812 672 1824 684
rect 1836 672 1848 684
rect 1860 672 1872 684
rect 1884 672 1896 684
rect 1908 672 1920 684
rect 1932 672 1944 684
rect 1956 672 1968 684
rect 1980 672 1992 684
rect 2004 672 2016 684
rect 2028 672 2040 684
rect 2052 672 2064 684
rect 2076 672 2088 684
rect 2100 672 2112 684
rect 2124 672 2136 684
rect 2148 672 2160 684
rect 2172 672 2184 684
rect 2196 672 2208 684
rect 2220 672 2232 684
rect 2244 672 2256 684
rect 2268 672 2280 684
rect 2292 672 2304 684
rect 2316 672 2328 684
rect 2340 672 2352 684
rect 2364 672 2376 684
rect 2388 672 2400 684
rect 2412 672 2424 684
rect 2436 672 2448 684
rect 2460 672 2472 684
rect 2484 672 2496 684
rect 2508 672 2520 684
rect 2532 672 2544 684
rect 2556 672 2568 684
rect 2580 672 2592 684
rect 2604 672 2616 684
rect 2628 672 2640 684
rect 2652 672 2664 684
rect 2676 672 2688 684
rect 2700 672 2712 684
rect 2724 672 2736 684
rect 2748 672 2760 684
rect 2772 672 2784 684
rect 2796 672 2808 684
rect 2820 672 2832 684
rect 2844 672 2856 684
rect 2868 672 2880 684
rect 2892 672 2904 684
rect 2916 672 2928 684
rect 2940 672 2952 684
rect -996 -264 -984 -252
rect -972 -264 -960 -252
rect -948 -264 -936 -252
rect -924 -264 -912 -252
rect -900 -264 -888 -252
rect -876 -264 -864 -252
rect -852 -264 -840 -252
rect -828 -264 -816 -252
rect -804 -264 -792 -252
rect -780 -264 -768 -252
rect -756 -264 -744 -252
rect -732 -264 -720 -252
rect -708 -264 -696 -252
rect -684 -264 -672 -252
rect -660 -264 -648 -252
rect -636 -264 -624 -252
rect -612 -264 -600 -252
rect -588 -264 -576 -252
rect -564 -264 -552 -252
rect -540 -264 -528 -252
rect -516 -264 -504 -252
rect -492 -264 -480 -252
rect -468 -264 -456 -252
rect -444 -264 -432 -252
rect -420 -264 -408 -252
rect -396 -264 -384 -252
rect -372 -264 -360 -252
rect -348 -264 -336 -252
rect -324 -264 -312 -252
rect -300 -264 -288 -252
rect -276 -264 -264 -252
rect -252 -264 -240 -252
rect -228 -264 -216 -252
rect -204 -264 -192 -252
rect -180 -264 -168 -252
rect -156 -264 -144 -252
rect -132 -264 -120 -252
rect -108 -264 -96 -252
rect -84 -264 -72 -252
rect -60 -264 -48 -252
rect -36 -264 -24 -252
rect -12 -264 0 -252
rect 12 -264 24 -252
rect 36 -264 48 -252
rect 60 -264 72 -252
rect 84 -264 96 -252
rect 108 -264 120 -252
rect 132 -264 144 -252
rect 156 -264 168 -252
rect 180 -264 192 -252
rect 204 -264 216 -252
rect 228 -264 240 -252
rect 252 -264 264 -252
rect 276 -264 288 -252
rect 300 -264 312 -252
rect 324 -264 336 -252
rect 348 -264 360 -252
rect 372 -264 384 -252
rect 396 -264 408 -252
rect 420 -264 432 -252
rect 444 -264 456 -252
rect 468 -264 480 -252
rect 492 -264 504 -252
rect 516 -264 528 -252
rect 540 -264 552 -252
rect 564 -264 576 -252
rect 588 -264 600 -252
rect 612 -264 624 -252
rect 636 -264 648 -252
rect 660 -264 672 -252
rect 684 -264 696 -252
rect 708 -264 720 -252
rect 732 -264 744 -252
rect 756 -264 768 -252
rect 780 -264 792 -252
rect 804 -264 816 -252
rect 828 -264 840 -252
rect 852 -264 864 -252
rect 876 -264 888 -252
rect 900 -264 912 -252
rect 924 -264 936 -252
rect 948 -264 960 -252
rect 972 -264 984 -252
rect 996 -264 1008 -252
rect 1020 -264 1032 -252
rect 1044 -264 1056 -252
rect 1068 -264 1080 -252
rect 1092 -264 1104 -252
rect 1116 -264 1128 -252
rect 1140 -264 1152 -252
rect 1164 -264 1176 -252
rect 1188 -264 1200 -252
rect 1212 -264 1224 -252
rect 1236 -264 1248 -252
rect 1260 -264 1272 -252
rect 1284 -264 1296 -252
rect 1308 -264 1320 -252
rect 1332 -264 1344 -252
rect 1356 -264 1368 -252
rect 1380 -264 1392 -252
rect 1404 -264 1416 -252
rect 1428 -264 1440 -252
rect 1452 -264 1464 -252
rect 1476 -264 1488 -252
rect 1500 -264 1512 -252
rect 1524 -264 1536 -252
rect 1548 -264 1560 -252
rect 1572 -264 1584 -252
rect 1596 -264 1608 -252
rect 1620 -264 1632 -252
rect 1644 -264 1656 -252
rect 1668 -264 1680 -252
rect 1692 -264 1704 -252
rect 1716 -264 1728 -252
rect 1740 -264 1752 -252
rect 1764 -264 1776 -252
rect 1788 -264 1800 -252
rect 1812 -264 1824 -252
rect 1836 -264 1848 -252
rect 1860 -264 1872 -252
rect 1884 -264 1896 -252
rect 1908 -264 1920 -252
rect 1932 -264 1944 -252
rect 1956 -264 1968 -252
rect 1980 -264 1992 -252
rect 2004 -264 2016 -252
rect 2028 -264 2040 -252
rect 2052 -264 2064 -252
rect 2076 -264 2088 -252
rect 2100 -264 2112 -252
rect 2124 -264 2136 -252
rect 2148 -264 2160 -252
rect 2172 -264 2184 -252
rect 2196 -264 2208 -252
rect 2220 -264 2232 -252
rect 2244 -264 2256 -252
rect 2268 -264 2280 -252
rect 2292 -264 2304 -252
rect 2316 -264 2328 -252
rect 2340 -264 2352 -252
rect 2364 -264 2376 -252
rect 2388 -264 2400 -252
rect 2412 -264 2424 -252
rect 2436 -264 2448 -252
rect 2460 -264 2472 -252
rect 2484 -264 2496 -252
rect 2508 -264 2520 -252
rect 2532 -264 2544 -252
rect 2556 -264 2568 -252
rect 2580 -264 2592 -252
rect 2604 -264 2616 -252
rect 2628 -264 2640 -252
rect 2652 -264 2664 -252
rect 2676 -264 2688 -252
rect 2700 -264 2712 -252
rect 2724 -264 2736 -252
rect 2748 -264 2760 -252
rect 2772 -264 2784 -252
rect 2796 -264 2808 -252
rect 2820 -264 2832 -252
rect 2844 -264 2856 -252
rect 2868 -264 2880 -252
rect 2892 -264 2904 -252
rect 2916 -264 2928 -252
rect 2940 -264 2952 -252
rect -996 -300 -984 -288
rect -972 -300 -960 -288
rect -948 -300 -936 -288
rect -924 -300 -912 -288
rect -900 -300 -888 -288
rect -876 -300 -864 -288
rect -852 -300 -840 -288
rect -828 -300 -816 -288
rect -804 -300 -792 -288
rect -780 -300 -768 -288
rect -756 -300 -744 -288
rect -732 -300 -720 -288
rect -708 -300 -696 -288
rect -684 -300 -672 -288
rect -660 -300 -648 -288
rect -636 -300 -624 -288
rect -612 -300 -600 -288
rect -588 -300 -576 -288
rect -564 -300 -552 -288
rect -540 -300 -528 -288
rect -516 -300 -504 -288
rect -492 -300 -480 -288
rect -468 -300 -456 -288
rect -444 -300 -432 -288
rect -420 -300 -408 -288
rect -396 -300 -384 -288
rect -372 -300 -360 -288
rect -348 -300 -336 -288
rect -324 -300 -312 -288
rect -300 -300 -288 -288
rect -276 -300 -264 -288
rect -252 -300 -240 -288
rect -228 -300 -216 -288
rect -204 -300 -192 -288
rect -180 -300 -168 -288
rect -156 -300 -144 -288
rect -132 -300 -120 -288
rect -108 -300 -96 -288
rect -84 -300 -72 -288
rect -60 -300 -48 -288
rect -36 -300 -24 -288
rect -12 -300 0 -288
rect 12 -300 24 -288
rect 36 -300 48 -288
rect 60 -300 72 -288
rect 84 -300 96 -288
rect 108 -300 120 -288
rect 132 -300 144 -288
rect 156 -300 168 -288
rect 180 -300 192 -288
rect 204 -300 216 -288
rect 228 -300 240 -288
rect 252 -300 264 -288
rect 276 -300 288 -288
rect 300 -300 312 -288
rect 324 -300 336 -288
rect 348 -300 360 -288
rect 372 -300 384 -288
rect 396 -300 408 -288
rect 420 -300 432 -288
rect 444 -300 456 -288
rect 468 -300 480 -288
rect 492 -300 504 -288
rect 516 -300 528 -288
rect 540 -300 552 -288
rect 564 -300 576 -288
rect 588 -300 600 -288
rect 612 -300 624 -288
rect 636 -300 648 -288
rect 660 -300 672 -288
rect 684 -300 696 -288
rect 708 -300 720 -288
rect 732 -300 744 -288
rect 756 -300 768 -288
rect 780 -300 792 -288
rect 804 -300 816 -288
rect 828 -300 840 -288
rect 852 -300 864 -288
rect 876 -300 888 -288
rect 900 -300 912 -288
rect 924 -300 936 -288
rect 948 -300 960 -288
rect 972 -300 984 -288
rect 996 -300 1008 -288
rect 1020 -300 1032 -288
rect 1044 -300 1056 -288
rect 1068 -300 1080 -288
rect 1092 -300 1104 -288
rect 1116 -300 1128 -288
rect 1140 -300 1152 -288
rect 1164 -300 1176 -288
rect 1188 -300 1200 -288
rect 1212 -300 1224 -288
rect 1236 -300 1248 -288
rect 1260 -300 1272 -288
rect 1284 -300 1296 -288
rect 1308 -300 1320 -288
rect 1332 -300 1344 -288
rect 1356 -300 1368 -288
rect 1380 -300 1392 -288
rect 1404 -300 1416 -288
rect 1428 -300 1440 -288
rect 1452 -300 1464 -288
rect 1476 -300 1488 -288
rect 1500 -300 1512 -288
rect 1524 -300 1536 -288
rect 1548 -300 1560 -288
rect 1572 -300 1584 -288
rect 1596 -300 1608 -288
rect 1620 -300 1632 -288
rect 1644 -300 1656 -288
rect 1668 -300 1680 -288
rect 1692 -300 1704 -288
rect 1716 -300 1728 -288
rect 1740 -300 1752 -288
rect 1764 -300 1776 -288
rect 1788 -300 1800 -288
rect 1812 -300 1824 -288
rect 1836 -300 1848 -288
rect 1860 -300 1872 -288
rect 1884 -300 1896 -288
rect 1908 -300 1920 -288
rect 1932 -300 1944 -288
rect 1956 -300 1968 -288
rect 1980 -300 1992 -288
rect 2004 -300 2016 -288
rect 2028 -300 2040 -288
rect 2052 -300 2064 -288
rect 2076 -300 2088 -288
rect 2100 -300 2112 -288
rect 2124 -300 2136 -288
rect 2148 -300 2160 -288
rect 2172 -300 2184 -288
rect 2196 -300 2208 -288
rect 2220 -300 2232 -288
rect 2244 -300 2256 -288
rect 2268 -300 2280 -288
rect 2292 -300 2304 -288
rect 2316 -300 2328 -288
rect 2340 -300 2352 -288
rect 2364 -300 2376 -288
rect 2388 -300 2400 -288
rect 2412 -300 2424 -288
rect 2436 -300 2448 -288
rect 2460 -300 2472 -288
rect 2484 -300 2496 -288
rect 2508 -300 2520 -288
rect 2532 -300 2544 -288
rect 2556 -300 2568 -288
rect 2580 -300 2592 -288
rect 2604 -300 2616 -288
rect 2628 -300 2640 -288
rect 2652 -300 2664 -288
rect 2676 -300 2688 -288
rect 2700 -300 2712 -288
rect 2724 -300 2736 -288
rect 2748 -300 2760 -288
rect 2772 -300 2784 -288
rect 2796 -300 2808 -288
rect 2820 -300 2832 -288
rect 2844 -300 2856 -288
rect 2868 -300 2880 -288
rect 2892 -300 2904 -288
rect 2916 -300 2928 -288
rect 2940 -300 2952 -288
rect -996 -336 -984 -324
rect -972 -336 -960 -324
rect -948 -336 -936 -324
rect -924 -336 -912 -324
rect -900 -336 -888 -324
rect -876 -336 -864 -324
rect -852 -336 -840 -324
rect -828 -336 -816 -324
rect -804 -336 -792 -324
rect -780 -336 -768 -324
rect -756 -336 -744 -324
rect -732 -336 -720 -324
rect -708 -336 -696 -324
rect -684 -336 -672 -324
rect -660 -336 -648 -324
rect -636 -336 -624 -324
rect -612 -336 -600 -324
rect -588 -336 -576 -324
rect -564 -336 -552 -324
rect -540 -336 -528 -324
rect -516 -336 -504 -324
rect -492 -336 -480 -324
rect -468 -336 -456 -324
rect -444 -336 -432 -324
rect -420 -336 -408 -324
rect -396 -336 -384 -324
rect -372 -336 -360 -324
rect -348 -336 -336 -324
rect -324 -336 -312 -324
rect -300 -336 -288 -324
rect -276 -336 -264 -324
rect -252 -336 -240 -324
rect -228 -336 -216 -324
rect -204 -336 -192 -324
rect -180 -336 -168 -324
rect -156 -336 -144 -324
rect -132 -336 -120 -324
rect -108 -336 -96 -324
rect -84 -336 -72 -324
rect -60 -336 -48 -324
rect -36 -336 -24 -324
rect -12 -336 0 -324
rect 12 -336 24 -324
rect 36 -336 48 -324
rect 60 -336 72 -324
rect 84 -336 96 -324
rect 108 -336 120 -324
rect 132 -336 144 -324
rect 156 -336 168 -324
rect 180 -336 192 -324
rect 204 -336 216 -324
rect 228 -336 240 -324
rect 252 -336 264 -324
rect 276 -336 288 -324
rect 300 -336 312 -324
rect 324 -336 336 -324
rect 348 -336 360 -324
rect 372 -336 384 -324
rect 396 -336 408 -324
rect 420 -336 432 -324
rect 444 -336 456 -324
rect 468 -336 480 -324
rect 492 -336 504 -324
rect 516 -336 528 -324
rect 540 -336 552 -324
rect 564 -336 576 -324
rect 588 -336 600 -324
rect 612 -336 624 -324
rect 636 -336 648 -324
rect 660 -336 672 -324
rect 684 -336 696 -324
rect 708 -336 720 -324
rect 732 -336 744 -324
rect 756 -336 768 -324
rect 780 -336 792 -324
rect 804 -336 816 -324
rect 828 -336 840 -324
rect 852 -336 864 -324
rect 876 -336 888 -324
rect 900 -336 912 -324
rect 924 -336 936 -324
rect 948 -336 960 -324
rect 972 -336 984 -324
rect 996 -336 1008 -324
rect 1020 -336 1032 -324
rect 1044 -336 1056 -324
rect 1068 -336 1080 -324
rect 1092 -336 1104 -324
rect 1116 -336 1128 -324
rect 1140 -336 1152 -324
rect 1164 -336 1176 -324
rect 1188 -336 1200 -324
rect 1212 -336 1224 -324
rect 1236 -336 1248 -324
rect 1260 -336 1272 -324
rect 1284 -336 1296 -324
rect 1308 -336 1320 -324
rect 1332 -336 1344 -324
rect 1356 -336 1368 -324
rect 1380 -336 1392 -324
rect 1404 -336 1416 -324
rect 1428 -336 1440 -324
rect 1452 -336 1464 -324
rect 1476 -336 1488 -324
rect 1500 -336 1512 -324
rect 1524 -336 1536 -324
rect 1548 -336 1560 -324
rect 1572 -336 1584 -324
rect 1596 -336 1608 -324
rect 1620 -336 1632 -324
rect 1644 -336 1656 -324
rect 1668 -336 1680 -324
rect 1692 -336 1704 -324
rect 1716 -336 1728 -324
rect 1740 -336 1752 -324
rect 1764 -336 1776 -324
rect 1788 -336 1800 -324
rect 1812 -336 1824 -324
rect 1836 -336 1848 -324
rect 1860 -336 1872 -324
rect 1884 -336 1896 -324
rect 1908 -336 1920 -324
rect 1932 -336 1944 -324
rect 1956 -336 1968 -324
rect 1980 -336 1992 -324
rect 2004 -336 2016 -324
rect 2028 -336 2040 -324
rect 2052 -336 2064 -324
rect 2076 -336 2088 -324
rect 2100 -336 2112 -324
rect 2124 -336 2136 -324
rect 2148 -336 2160 -324
rect 2172 -336 2184 -324
rect 2196 -336 2208 -324
rect 2220 -336 2232 -324
rect 2244 -336 2256 -324
rect 2268 -336 2280 -324
rect 2292 -336 2304 -324
rect 2316 -336 2328 -324
rect 2340 -336 2352 -324
rect 2364 -336 2376 -324
rect 2388 -336 2400 -324
rect 2412 -336 2424 -324
rect 2436 -336 2448 -324
rect 2460 -336 2472 -324
rect 2484 -336 2496 -324
rect 2508 -336 2520 -324
rect 2532 -336 2544 -324
rect 2556 -336 2568 -324
rect 2580 -336 2592 -324
rect 2604 -336 2616 -324
rect 2628 -336 2640 -324
rect 2652 -336 2664 -324
rect 2676 -336 2688 -324
rect 2700 -336 2712 -324
rect 2724 -336 2736 -324
rect 2748 -336 2760 -324
rect 2772 -336 2784 -324
rect 2796 -336 2808 -324
rect 2820 -336 2832 -324
rect 2844 -336 2856 -324
rect 2868 -336 2880 -324
rect 2892 -336 2904 -324
rect 2916 -336 2928 -324
rect 2940 -336 2952 -324
rect -996 -372 -984 -360
rect -972 -372 -960 -360
rect -948 -372 -936 -360
rect -924 -372 -912 -360
rect -900 -372 -888 -360
rect -876 -372 -864 -360
rect -852 -372 -840 -360
rect -828 -372 -816 -360
rect -804 -372 -792 -360
rect -780 -372 -768 -360
rect -756 -372 -744 -360
rect -732 -372 -720 -360
rect -708 -372 -696 -360
rect -684 -372 -672 -360
rect -660 -372 -648 -360
rect -636 -372 -624 -360
rect -612 -372 -600 -360
rect -588 -372 -576 -360
rect -564 -372 -552 -360
rect -540 -372 -528 -360
rect -516 -372 -504 -360
rect -492 -372 -480 -360
rect -468 -372 -456 -360
rect -444 -372 -432 -360
rect -420 -372 -408 -360
rect -396 -372 -384 -360
rect -372 -372 -360 -360
rect -348 -372 -336 -360
rect -324 -372 -312 -360
rect -300 -372 -288 -360
rect -276 -372 -264 -360
rect -252 -372 -240 -360
rect -228 -372 -216 -360
rect -204 -372 -192 -360
rect -180 -372 -168 -360
rect -156 -372 -144 -360
rect -132 -372 -120 -360
rect -108 -372 -96 -360
rect -84 -372 -72 -360
rect -60 -372 -48 -360
rect -36 -372 -24 -360
rect -12 -372 0 -360
rect 12 -372 24 -360
rect 36 -372 48 -360
rect 60 -372 72 -360
rect 84 -372 96 -360
rect 108 -372 120 -360
rect 132 -372 144 -360
rect 156 -372 168 -360
rect 180 -372 192 -360
rect 204 -372 216 -360
rect 228 -372 240 -360
rect 252 -372 264 -360
rect 276 -372 288 -360
rect 300 -372 312 -360
rect 324 -372 336 -360
rect 348 -372 360 -360
rect 372 -372 384 -360
rect 396 -372 408 -360
rect 420 -372 432 -360
rect 444 -372 456 -360
rect 468 -372 480 -360
rect 492 -372 504 -360
rect 516 -372 528 -360
rect 540 -372 552 -360
rect 564 -372 576 -360
rect 588 -372 600 -360
rect 612 -372 624 -360
rect 636 -372 648 -360
rect 660 -372 672 -360
rect 684 -372 696 -360
rect 708 -372 720 -360
rect 732 -372 744 -360
rect 756 -372 768 -360
rect 780 -372 792 -360
rect 804 -372 816 -360
rect 828 -372 840 -360
rect 852 -372 864 -360
rect 876 -372 888 -360
rect 900 -372 912 -360
rect 924 -372 936 -360
rect 948 -372 960 -360
rect 972 -372 984 -360
rect 996 -372 1008 -360
rect 1020 -372 1032 -360
rect 1044 -372 1056 -360
rect 1068 -372 1080 -360
rect 1092 -372 1104 -360
rect 1116 -372 1128 -360
rect 1140 -372 1152 -360
rect 1164 -372 1176 -360
rect 1188 -372 1200 -360
rect 1212 -372 1224 -360
rect 1236 -372 1248 -360
rect 1260 -372 1272 -360
rect 1284 -372 1296 -360
rect 1308 -372 1320 -360
rect 1332 -372 1344 -360
rect 1356 -372 1368 -360
rect 1380 -372 1392 -360
rect 1404 -372 1416 -360
rect 1428 -372 1440 -360
rect 1452 -372 1464 -360
rect 1476 -372 1488 -360
rect 1500 -372 1512 -360
rect 1524 -372 1536 -360
rect 1548 -372 1560 -360
rect 1572 -372 1584 -360
rect 1596 -372 1608 -360
rect 1620 -372 1632 -360
rect 1644 -372 1656 -360
rect 1668 -372 1680 -360
rect 1692 -372 1704 -360
rect 1716 -372 1728 -360
rect 1740 -372 1752 -360
rect 1764 -372 1776 -360
rect 1788 -372 1800 -360
rect 1812 -372 1824 -360
rect 1836 -372 1848 -360
rect 1860 -372 1872 -360
rect 1884 -372 1896 -360
rect 1908 -372 1920 -360
rect 1932 -372 1944 -360
rect 1956 -372 1968 -360
rect 1980 -372 1992 -360
rect 2004 -372 2016 -360
rect 2028 -372 2040 -360
rect 2052 -372 2064 -360
rect 2076 -372 2088 -360
rect 2100 -372 2112 -360
rect 2124 -372 2136 -360
rect 2148 -372 2160 -360
rect 2172 -372 2184 -360
rect 2196 -372 2208 -360
rect 2220 -372 2232 -360
rect 2244 -372 2256 -360
rect 2268 -372 2280 -360
rect 2292 -372 2304 -360
rect 2316 -372 2328 -360
rect 2340 -372 2352 -360
rect 2364 -372 2376 -360
rect 2388 -372 2400 -360
rect 2412 -372 2424 -360
rect 2436 -372 2448 -360
rect 2460 -372 2472 -360
rect 2484 -372 2496 -360
rect 2508 -372 2520 -360
rect 2532 -372 2544 -360
rect 2556 -372 2568 -360
rect 2580 -372 2592 -360
rect 2604 -372 2616 -360
rect 2628 -372 2640 -360
rect 2652 -372 2664 -360
rect 2676 -372 2688 -360
rect 2700 -372 2712 -360
rect 2724 -372 2736 -360
rect 2748 -372 2760 -360
rect 2772 -372 2784 -360
rect 2796 -372 2808 -360
rect 2820 -372 2832 -360
rect 2844 -372 2856 -360
rect 2868 -372 2880 -360
rect 2892 -372 2904 -360
rect 2916 -372 2928 -360
rect 2940 -372 2952 -360
<< metal3 >>
rect -1044 492 -1032 552
rect -1044 438 -1032 456
rect -1044 420 -1032 432
rect -1044 288 -1032 300
rect -1104 250 -1032 252
rect -1104 224 -1102 250
rect -1094 224 -1054 250
rect -1046 224 -1032 250
rect -1104 222 -1032 224
rect -1104 214 -1032 216
rect -1104 206 -1078 214
rect -1070 206 -1032 214
rect -1104 204 -1032 206
rect -1104 196 -1032 198
rect -1104 170 -1102 196
rect -1094 170 -1054 196
rect -1046 170 -1032 196
rect -1104 168 -1032 170
rect -1044 120 -1032 132
rect -1044 72 -1032 84
rect -1104 34 -1032 36
rect -1104 8 -1102 34
rect -1094 8 -1054 34
rect -1046 8 -1032 34
rect -1104 6 -1032 8
rect -1104 -2 -1032 0
rect -1104 -10 -1078 -2
rect -1070 -10 -1032 -2
rect -1104 -12 -1032 -10
rect -1104 -20 -1032 -18
rect -1104 -46 -1102 -20
rect -1094 -46 -1054 -20
rect -1046 -46 -1032 -20
rect -1104 -48 -1032 -46
rect -1044 -168 -1032 -108
<< via3 >>
rect -1102 224 -1094 250
rect -1054 224 -1046 250
rect -144 228 -132 252
rect -72 228 -60 252
rect 576 228 588 252
rect 648 228 660 252
rect 1296 228 1308 252
rect 1368 228 1380 252
rect 2016 228 2028 252
rect 2088 228 2100 252
rect -1078 206 -1070 214
rect -744 204 -732 216
rect -672 204 -660 216
rect -432 204 -420 216
rect 216 204 228 216
rect 288 204 300 216
rect 936 204 948 216
rect 1008 204 1020 216
rect 1656 204 1668 216
rect 1728 204 1740 216
rect 2376 204 2388 216
rect 2616 204 2628 216
rect 2688 204 2700 216
rect -1102 170 -1094 196
rect -1054 170 -1046 196
rect -144 168 -132 192
rect -72 168 -60 192
rect 576 168 588 192
rect 648 168 660 192
rect 1296 168 1308 192
rect 1368 168 1380 192
rect 2016 168 2028 192
rect 2088 168 2100 192
rect -912 120 -900 132
rect -864 120 -852 132
rect -384 120 -372 132
rect 168 120 180 132
rect 336 120 348 132
rect 888 120 900 132
rect 1056 120 1068 132
rect 1608 120 1620 132
rect 1776 120 1788 132
rect 2328 120 2340 132
rect 2808 120 2820 132
rect 2856 120 2868 132
rect -552 72 -540 84
rect -504 72 -492 84
rect -312 72 -300 84
rect 96 72 108 84
rect 408 72 420 84
rect 816 72 828 84
rect 1128 72 1140 84
rect 1536 72 1548 84
rect 1848 72 1860 84
rect 2256 72 2268 84
rect 2448 72 2460 84
rect 2496 72 2508 84
rect -1102 8 -1094 34
rect -1054 8 -1046 34
rect -192 12 -180 36
rect -24 12 -12 36
rect 528 12 540 36
rect 696 12 708 36
rect 1248 12 1260 36
rect 1416 12 1428 36
rect 1968 12 1980 36
rect 2136 12 2148 36
rect -1078 -10 -1070 -2
rect -792 -12 -780 0
rect -624 -12 -612 0
rect -264 -12 -252 0
rect 48 -12 60 0
rect 456 -12 468 0
rect 768 -12 780 0
rect 1176 -12 1188 0
rect 1488 -12 1500 0
rect 1896 -12 1908 0
rect 2208 -12 2220 0
rect 2568 -12 2580 0
rect 2736 -12 2748 0
rect -1102 -46 -1094 -20
rect -1054 -46 -1046 -20
rect -192 -48 -180 -24
rect -24 -48 -12 -24
rect 528 -48 540 -24
rect 696 -48 708 -24
rect 1248 -48 1260 -24
rect 1416 -48 1428 -24
rect 1968 -48 1980 -24
rect 2136 -48 2148 -24
<< metal4 >>
rect -1020 804 2988 816
rect -1104 660 -1092 672
rect -1104 612 -1092 648
rect -1104 250 -1092 600
rect -1104 224 -1102 250
rect -1094 224 -1092 250
rect -1104 196 -1092 224
rect -1104 170 -1102 196
rect -1094 170 -1092 196
rect -1104 168 -1092 170
rect -1080 636 -1068 672
rect -1080 214 -1068 624
rect -1080 206 -1078 214
rect -1070 206 -1068 214
rect -1080 168 -1068 206
rect -1056 660 -1044 672
rect -1056 612 -1044 648
rect -1020 660 -1008 804
rect 2976 660 2988 804
rect -1020 636 2988 660
rect -1020 624 -1008 636
rect -996 624 -984 636
rect -972 624 -960 636
rect -948 624 -936 636
rect -924 624 -912 636
rect -900 624 -888 636
rect -876 624 -864 636
rect -852 624 -840 636
rect -828 624 -804 636
rect -792 624 -780 636
rect -768 624 -756 636
rect -744 624 -732 636
rect -720 624 -708 636
rect -696 624 -684 636
rect -672 624 -660 636
rect -648 624 -636 636
rect -624 624 -612 636
rect -600 624 -588 636
rect -576 624 -564 636
rect -552 624 -540 636
rect -528 624 -516 636
rect -504 624 -492 636
rect -480 624 -468 636
rect -456 624 -444 636
rect -432 624 -408 636
rect -396 624 -384 636
rect -372 624 -360 636
rect -348 624 -336 636
rect -324 624 -312 636
rect -300 624 -288 636
rect -276 624 -264 636
rect -252 624 -240 636
rect -228 624 -204 636
rect -192 624 -180 636
rect -168 624 -156 636
rect -144 624 -132 636
rect -120 624 -108 636
rect -96 624 -84 636
rect -72 624 -60 636
rect -48 624 -36 636
rect -24 624 -12 636
rect 0 624 12 636
rect 24 624 36 636
rect 48 624 60 636
rect 72 624 84 636
rect 96 624 108 636
rect 120 624 132 636
rect 144 624 156 636
rect 168 624 180 636
rect 192 624 204 636
rect 216 624 228 636
rect 240 624 252 636
rect 264 624 276 636
rect 288 624 300 636
rect 312 624 324 636
rect 336 624 348 636
rect 360 624 384 636
rect 396 624 408 636
rect 420 624 432 636
rect 444 624 456 636
rect 468 624 480 636
rect 492 624 504 636
rect 516 624 528 636
rect 540 624 552 636
rect 564 624 576 636
rect 588 624 600 636
rect 612 624 624 636
rect 636 624 648 636
rect 660 624 672 636
rect 684 624 696 636
rect 708 624 720 636
rect 732 624 744 636
rect 756 624 768 636
rect 780 624 792 636
rect 804 624 816 636
rect 828 624 840 636
rect 852 624 864 636
rect 876 624 888 636
rect 900 624 912 636
rect 924 624 936 636
rect 948 624 972 636
rect 984 624 996 636
rect 1008 624 1020 636
rect 1032 624 1044 636
rect 1056 624 1068 636
rect 1080 624 1092 636
rect 1104 624 1116 636
rect 1128 624 1140 636
rect 1152 624 1164 636
rect 1176 624 1188 636
rect 1200 624 1212 636
rect 1224 624 1236 636
rect 1248 624 1260 636
rect 1272 624 1284 636
rect 1296 624 1308 636
rect 1320 624 1332 636
rect 1344 624 1356 636
rect 1368 624 1380 636
rect 1392 624 1404 636
rect 1416 624 1428 636
rect 1440 624 1452 636
rect 1464 624 1476 636
rect 1488 624 1500 636
rect 1512 624 1524 636
rect 1536 624 1560 636
rect 1572 624 1584 636
rect 1596 624 1608 636
rect 1620 624 1632 636
rect 1644 624 1656 636
rect 1668 624 1680 636
rect 1692 624 1704 636
rect 1716 624 1728 636
rect 1740 624 1752 636
rect 1764 624 1776 636
rect 1788 624 1800 636
rect 1812 624 1824 636
rect 1836 624 1848 636
rect 1860 624 1872 636
rect 1884 624 1896 636
rect 1908 624 1920 636
rect 1932 624 1956 636
rect 1968 624 1980 636
rect 1992 624 2004 636
rect 2016 624 2028 636
rect 2040 624 2052 636
rect 2064 624 2076 636
rect 2088 624 2100 636
rect 2112 624 2124 636
rect 2136 624 2160 636
rect 2172 624 2184 636
rect 2196 624 2208 636
rect 2220 624 2232 636
rect 2244 624 2256 636
rect 2268 624 2280 636
rect 2292 624 2304 636
rect 2316 624 2328 636
rect 2340 624 2352 636
rect 2364 624 2376 636
rect 2388 624 2400 636
rect 2412 624 2424 636
rect 2436 624 2448 636
rect 2460 624 2472 636
rect 2484 624 2496 636
rect 2508 624 2520 636
rect 2532 624 2544 636
rect 2556 624 2568 636
rect 2580 624 2592 636
rect 2604 624 2616 636
rect 2628 624 2640 636
rect 2652 624 2664 636
rect 2676 624 2688 636
rect 2700 624 2712 636
rect 2724 624 2748 636
rect 2760 624 2772 636
rect 2784 624 2796 636
rect 2808 624 2820 636
rect 2832 624 2844 636
rect 2856 624 2868 636
rect 2880 624 2892 636
rect 2904 624 2916 636
rect 2928 624 2940 636
rect 2952 624 2964 636
rect 2976 624 2988 636
rect -1020 612 2988 624
rect -1056 250 -1044 600
rect -1056 224 -1054 250
rect -1046 224 -1044 250
rect -1056 196 -1044 224
rect -1056 170 -1054 196
rect -1046 170 -1044 196
rect -1056 168 -1044 170
rect -1104 34 -1092 36
rect -1104 8 -1102 34
rect -1094 8 -1092 34
rect -1104 -20 -1092 8
rect -1104 -46 -1102 -20
rect -1094 -46 -1092 -20
rect -1104 -180 -1092 -46
rect -1104 -228 -1092 -192
rect -1104 -252 -1092 -240
rect -1080 -2 -1068 36
rect -1080 -10 -1078 -2
rect -1070 -10 -1068 -2
rect -1080 -204 -1068 -10
rect -1080 -252 -1068 -216
rect -1056 34 -1044 36
rect -1056 8 -1054 34
rect -1046 8 -1044 34
rect -1056 -20 -1044 8
rect -1056 -46 -1054 -20
rect -1046 -46 -1044 -20
rect -1056 -180 -1044 -46
rect -1056 -228 -1044 -192
rect -1056 -252 -1044 -240
rect -1020 -204 2988 -192
rect -1020 -216 -1008 -204
rect -996 -216 -984 -204
rect -972 -216 -960 -204
rect -948 -216 -936 -204
rect -924 -216 -912 -204
rect -900 -216 -888 -204
rect -876 -216 -864 -204
rect -852 -216 -840 -204
rect -828 -216 -804 -204
rect -792 -216 -780 -204
rect -768 -216 -756 -204
rect -744 -216 -732 -204
rect -720 -216 -708 -204
rect -696 -216 -684 -204
rect -672 -216 -660 -204
rect -648 -216 -636 -204
rect -624 -216 -612 -204
rect -600 -216 -588 -204
rect -576 -216 -564 -204
rect -552 -216 -540 -204
rect -528 -216 -516 -204
rect -504 -216 -492 -204
rect -480 -216 -468 -204
rect -456 -216 -444 -204
rect -432 -216 -408 -204
rect -396 -216 -384 -204
rect -372 -216 -360 -204
rect -348 -216 -336 -204
rect -324 -216 -312 -204
rect -300 -216 -288 -204
rect -276 -216 -264 -204
rect -252 -216 -240 -204
rect -228 -216 -204 -204
rect -192 -216 -180 -204
rect -168 -216 -156 -204
rect -144 -216 -132 -204
rect -120 -216 -108 -204
rect -96 -216 -84 -204
rect -72 -216 -60 -204
rect -48 -216 -36 -204
rect -24 -216 -12 -204
rect 0 -216 12 -204
rect 24 -216 36 -204
rect 48 -216 60 -204
rect 72 -216 84 -204
rect 96 -216 108 -204
rect 120 -216 132 -204
rect 144 -216 156 -204
rect 168 -216 180 -204
rect 192 -216 204 -204
rect 216 -216 228 -204
rect 240 -216 252 -204
rect 264 -216 276 -204
rect 288 -216 300 -204
rect 312 -216 324 -204
rect 336 -216 348 -204
rect 360 -216 384 -204
rect 396 -216 408 -204
rect 420 -216 432 -204
rect 444 -216 456 -204
rect 468 -216 480 -204
rect 492 -216 504 -204
rect 516 -216 528 -204
rect 540 -216 552 -204
rect 564 -216 576 -204
rect 588 -216 600 -204
rect 612 -216 624 -204
rect 636 -216 648 -204
rect 660 -216 672 -204
rect 684 -216 696 -204
rect 708 -216 720 -204
rect 732 -216 744 -204
rect 756 -216 768 -204
rect 780 -216 792 -204
rect 804 -216 816 -204
rect 828 -216 840 -204
rect 852 -216 864 -204
rect 876 -216 888 -204
rect 900 -216 912 -204
rect 924 -216 936 -204
rect 948 -216 972 -204
rect 984 -216 996 -204
rect 1008 -216 1020 -204
rect 1032 -216 1044 -204
rect 1056 -216 1068 -204
rect 1080 -216 1092 -204
rect 1104 -216 1116 -204
rect 1128 -216 1140 -204
rect 1152 -216 1164 -204
rect 1176 -216 1188 -204
rect 1200 -216 1212 -204
rect 1224 -216 1236 -204
rect 1248 -216 1260 -204
rect 1272 -216 1284 -204
rect 1296 -216 1308 -204
rect 1320 -216 1332 -204
rect 1344 -216 1356 -204
rect 1368 -216 1380 -204
rect 1392 -216 1404 -204
rect 1416 -216 1428 -204
rect 1440 -216 1452 -204
rect 1464 -216 1476 -204
rect 1488 -216 1500 -204
rect 1512 -216 1524 -204
rect 1536 -216 1560 -204
rect 1572 -216 1584 -204
rect 1596 -216 1608 -204
rect 1620 -216 1632 -204
rect 1644 -216 1656 -204
rect 1668 -216 1680 -204
rect 1692 -216 1704 -204
rect 1716 -216 1728 -204
rect 1740 -216 1752 -204
rect 1764 -216 1776 -204
rect 1788 -216 1800 -204
rect 1812 -216 1824 -204
rect 1836 -216 1848 -204
rect 1860 -216 1872 -204
rect 1884 -216 1896 -204
rect 1908 -216 1920 -204
rect 1932 -216 1956 -204
rect 1968 -216 1980 -204
rect 1992 -216 2004 -204
rect 2016 -216 2028 -204
rect 2040 -216 2052 -204
rect 2064 -216 2076 -204
rect 2088 -216 2100 -204
rect 2112 -216 2124 -204
rect 2136 -216 2160 -204
rect 2172 -216 2184 -204
rect 2196 -216 2208 -204
rect 2220 -216 2232 -204
rect 2244 -216 2256 -204
rect 2268 -216 2280 -204
rect 2292 -216 2304 -204
rect 2316 -216 2328 -204
rect 2340 -216 2352 -204
rect 2364 -216 2376 -204
rect 2388 -216 2400 -204
rect 2412 -216 2424 -204
rect 2436 -216 2448 -204
rect 2460 -216 2472 -204
rect 2484 -216 2496 -204
rect 2508 -216 2520 -204
rect 2532 -216 2544 -204
rect 2556 -216 2568 -204
rect 2580 -216 2592 -204
rect 2604 -216 2616 -204
rect 2628 -216 2640 -204
rect 2652 -216 2664 -204
rect 2676 -216 2688 -204
rect 2700 -216 2712 -204
rect 2724 -216 2748 -204
rect 2760 -216 2772 -204
rect 2784 -216 2796 -204
rect 2808 -216 2820 -204
rect 2832 -216 2844 -204
rect 2856 -216 2868 -204
rect 2880 -216 2892 -204
rect 2904 -216 2916 -204
rect 2928 -216 2940 -204
rect 2952 -216 2964 -204
rect 2976 -216 2988 -204
rect -1020 -240 2988 -216
rect -1020 -384 -1008 -240
rect 2976 -384 2988 -240
rect -1020 -396 2988 -384
<< via4 >>
rect -1104 648 -1092 660
rect -1104 600 -1092 612
rect -1080 624 -1068 636
rect -1056 648 -1044 660
rect -1008 624 -996 636
rect -984 624 -972 636
rect -960 624 -948 636
rect -936 624 -924 636
rect -912 624 -900 636
rect -888 624 -876 636
rect -864 624 -852 636
rect -840 624 -828 636
rect -804 624 -792 636
rect -780 624 -768 636
rect -756 624 -744 636
rect -732 624 -720 636
rect -708 624 -696 636
rect -684 624 -672 636
rect -660 624 -648 636
rect -636 624 -624 636
rect -612 624 -600 636
rect -588 624 -576 636
rect -564 624 -552 636
rect -540 624 -528 636
rect -516 624 -504 636
rect -492 624 -480 636
rect -468 624 -456 636
rect -444 624 -432 636
rect -408 624 -396 636
rect -384 624 -372 636
rect -360 624 -348 636
rect -336 624 -324 636
rect -312 624 -300 636
rect -288 624 -276 636
rect -264 624 -252 636
rect -240 624 -228 636
rect -204 624 -192 636
rect -180 624 -168 636
rect -156 624 -144 636
rect -132 624 -120 636
rect -108 624 -96 636
rect -84 624 -72 636
rect -60 624 -48 636
rect -36 624 -24 636
rect -12 624 0 636
rect 12 624 24 636
rect 36 624 48 636
rect 60 624 72 636
rect 84 624 96 636
rect 108 624 120 636
rect 132 624 144 636
rect 156 624 168 636
rect 180 624 192 636
rect 204 624 216 636
rect 228 624 240 636
rect 252 624 264 636
rect 276 624 288 636
rect 300 624 312 636
rect 324 624 336 636
rect 348 624 360 636
rect 384 624 396 636
rect 408 624 420 636
rect 432 624 444 636
rect 456 624 468 636
rect 480 624 492 636
rect 504 624 516 636
rect 528 624 540 636
rect 552 624 564 636
rect 576 624 588 636
rect 600 624 612 636
rect 624 624 636 636
rect 648 624 660 636
rect 672 624 684 636
rect 696 624 708 636
rect 720 624 732 636
rect 744 624 756 636
rect 768 624 780 636
rect 792 624 804 636
rect 816 624 828 636
rect 840 624 852 636
rect 864 624 876 636
rect 888 624 900 636
rect 912 624 924 636
rect 936 624 948 636
rect 972 624 984 636
rect 996 624 1008 636
rect 1020 624 1032 636
rect 1044 624 1056 636
rect 1068 624 1080 636
rect 1092 624 1104 636
rect 1116 624 1128 636
rect 1140 624 1152 636
rect 1164 624 1176 636
rect 1188 624 1200 636
rect 1212 624 1224 636
rect 1236 624 1248 636
rect 1260 624 1272 636
rect 1284 624 1296 636
rect 1308 624 1320 636
rect 1332 624 1344 636
rect 1356 624 1368 636
rect 1380 624 1392 636
rect 1404 624 1416 636
rect 1428 624 1440 636
rect 1452 624 1464 636
rect 1476 624 1488 636
rect 1500 624 1512 636
rect 1524 624 1536 636
rect 1560 624 1572 636
rect 1584 624 1596 636
rect 1608 624 1620 636
rect 1632 624 1644 636
rect 1656 624 1668 636
rect 1680 624 1692 636
rect 1704 624 1716 636
rect 1728 624 1740 636
rect 1752 624 1764 636
rect 1776 624 1788 636
rect 1800 624 1812 636
rect 1824 624 1836 636
rect 1848 624 1860 636
rect 1872 624 1884 636
rect 1896 624 1908 636
rect 1920 624 1932 636
rect 1956 624 1968 636
rect 1980 624 1992 636
rect 2004 624 2016 636
rect 2028 624 2040 636
rect 2052 624 2064 636
rect 2076 624 2088 636
rect 2100 624 2112 636
rect 2124 624 2136 636
rect 2160 624 2172 636
rect 2184 624 2196 636
rect 2208 624 2220 636
rect 2232 624 2244 636
rect 2256 624 2268 636
rect 2280 624 2292 636
rect 2304 624 2316 636
rect 2328 624 2340 636
rect 2352 624 2364 636
rect 2376 624 2388 636
rect 2400 624 2412 636
rect 2424 624 2436 636
rect 2448 624 2460 636
rect 2472 624 2484 636
rect 2496 624 2508 636
rect 2520 624 2532 636
rect 2544 624 2556 636
rect 2568 624 2580 636
rect 2592 624 2604 636
rect 2616 624 2628 636
rect 2640 624 2652 636
rect 2664 624 2676 636
rect 2688 624 2700 636
rect 2712 624 2724 636
rect 2748 624 2760 636
rect 2772 624 2784 636
rect 2796 624 2808 636
rect 2820 624 2832 636
rect 2844 624 2856 636
rect 2868 624 2880 636
rect 2892 624 2904 636
rect 2916 624 2928 636
rect 2940 624 2952 636
rect 2964 624 2976 636
rect -1056 600 -1044 612
rect -1104 -192 -1092 -180
rect -1104 -240 -1092 -228
rect -1080 -216 -1068 -204
rect -1056 -192 -1044 -180
rect -1056 -240 -1044 -228
rect -1008 -216 -996 -204
rect -984 -216 -972 -204
rect -960 -216 -948 -204
rect -936 -216 -924 -204
rect -912 -216 -900 -204
rect -888 -216 -876 -204
rect -864 -216 -852 -204
rect -840 -216 -828 -204
rect -804 -216 -792 -204
rect -780 -216 -768 -204
rect -756 -216 -744 -204
rect -732 -216 -720 -204
rect -708 -216 -696 -204
rect -684 -216 -672 -204
rect -660 -216 -648 -204
rect -636 -216 -624 -204
rect -612 -216 -600 -204
rect -588 -216 -576 -204
rect -564 -216 -552 -204
rect -540 -216 -528 -204
rect -516 -216 -504 -204
rect -492 -216 -480 -204
rect -468 -216 -456 -204
rect -444 -216 -432 -204
rect -408 -216 -396 -204
rect -384 -216 -372 -204
rect -360 -216 -348 -204
rect -336 -216 -324 -204
rect -312 -216 -300 -204
rect -288 -216 -276 -204
rect -264 -216 -252 -204
rect -240 -216 -228 -204
rect -204 -216 -192 -204
rect -180 -216 -168 -204
rect -156 -216 -144 -204
rect -132 -216 -120 -204
rect -108 -216 -96 -204
rect -84 -216 -72 -204
rect -60 -216 -48 -204
rect -36 -216 -24 -204
rect -12 -216 0 -204
rect 12 -216 24 -204
rect 36 -216 48 -204
rect 60 -216 72 -204
rect 84 -216 96 -204
rect 108 -216 120 -204
rect 132 -216 144 -204
rect 156 -216 168 -204
rect 180 -216 192 -204
rect 204 -216 216 -204
rect 228 -216 240 -204
rect 252 -216 264 -204
rect 276 -216 288 -204
rect 300 -216 312 -204
rect 324 -216 336 -204
rect 348 -216 360 -204
rect 384 -216 396 -204
rect 408 -216 420 -204
rect 432 -216 444 -204
rect 456 -216 468 -204
rect 480 -216 492 -204
rect 504 -216 516 -204
rect 528 -216 540 -204
rect 552 -216 564 -204
rect 576 -216 588 -204
rect 600 -216 612 -204
rect 624 -216 636 -204
rect 648 -216 660 -204
rect 672 -216 684 -204
rect 696 -216 708 -204
rect 720 -216 732 -204
rect 744 -216 756 -204
rect 768 -216 780 -204
rect 792 -216 804 -204
rect 816 -216 828 -204
rect 840 -216 852 -204
rect 864 -216 876 -204
rect 888 -216 900 -204
rect 912 -216 924 -204
rect 936 -216 948 -204
rect 972 -216 984 -204
rect 996 -216 1008 -204
rect 1020 -216 1032 -204
rect 1044 -216 1056 -204
rect 1068 -216 1080 -204
rect 1092 -216 1104 -204
rect 1116 -216 1128 -204
rect 1140 -216 1152 -204
rect 1164 -216 1176 -204
rect 1188 -216 1200 -204
rect 1212 -216 1224 -204
rect 1236 -216 1248 -204
rect 1260 -216 1272 -204
rect 1284 -216 1296 -204
rect 1308 -216 1320 -204
rect 1332 -216 1344 -204
rect 1356 -216 1368 -204
rect 1380 -216 1392 -204
rect 1404 -216 1416 -204
rect 1428 -216 1440 -204
rect 1452 -216 1464 -204
rect 1476 -216 1488 -204
rect 1500 -216 1512 -204
rect 1524 -216 1536 -204
rect 1560 -216 1572 -204
rect 1584 -216 1596 -204
rect 1608 -216 1620 -204
rect 1632 -216 1644 -204
rect 1656 -216 1668 -204
rect 1680 -216 1692 -204
rect 1704 -216 1716 -204
rect 1728 -216 1740 -204
rect 1752 -216 1764 -204
rect 1776 -216 1788 -204
rect 1800 -216 1812 -204
rect 1824 -216 1836 -204
rect 1848 -216 1860 -204
rect 1872 -216 1884 -204
rect 1896 -216 1908 -204
rect 1920 -216 1932 -204
rect 1956 -216 1968 -204
rect 1980 -216 1992 -204
rect 2004 -216 2016 -204
rect 2028 -216 2040 -204
rect 2052 -216 2064 -204
rect 2076 -216 2088 -204
rect 2100 -216 2112 -204
rect 2124 -216 2136 -204
rect 2160 -216 2172 -204
rect 2184 -216 2196 -204
rect 2208 -216 2220 -204
rect 2232 -216 2244 -204
rect 2256 -216 2268 -204
rect 2280 -216 2292 -204
rect 2304 -216 2316 -204
rect 2328 -216 2340 -204
rect 2352 -216 2364 -204
rect 2376 -216 2388 -204
rect 2400 -216 2412 -204
rect 2424 -216 2436 -204
rect 2448 -216 2460 -204
rect 2472 -216 2484 -204
rect 2496 -216 2508 -204
rect 2520 -216 2532 -204
rect 2544 -216 2556 -204
rect 2568 -216 2580 -204
rect 2592 -216 2604 -204
rect 2616 -216 2628 -204
rect 2640 -216 2652 -204
rect 2664 -216 2676 -204
rect 2688 -216 2700 -204
rect 2712 -216 2724 -204
rect 2748 -216 2760 -204
rect 2772 -216 2784 -204
rect 2796 -216 2808 -204
rect 2820 -216 2832 -204
rect 2844 -216 2856 -204
rect 2868 -216 2880 -204
rect 2892 -216 2904 -204
rect 2916 -216 2928 -204
rect 2940 -216 2952 -204
rect 2964 -216 2976 -204
<< metal5 >>
rect -1020 792 2988 816
rect -1020 780 -996 792
rect -984 780 -972 792
rect -960 780 -948 792
rect -936 780 -924 792
rect -912 780 -900 792
rect -888 780 -876 792
rect -864 780 -852 792
rect -840 780 -828 792
rect -816 780 -804 792
rect -792 780 -780 792
rect -768 780 -756 792
rect -744 780 -732 792
rect -720 780 -708 792
rect -696 780 -684 792
rect -672 780 -660 792
rect -648 780 -636 792
rect -624 780 -612 792
rect -600 780 -588 792
rect -576 780 -564 792
rect -552 780 -540 792
rect -528 780 -516 792
rect -504 780 -492 792
rect -480 780 -468 792
rect -456 780 -444 792
rect -432 780 -420 792
rect -408 780 -396 792
rect -384 780 -372 792
rect -360 780 -348 792
rect -336 780 -324 792
rect -312 780 -300 792
rect -288 780 -276 792
rect -264 780 -252 792
rect -240 780 -228 792
rect -216 780 -204 792
rect -192 780 -180 792
rect -168 780 -156 792
rect -144 780 -132 792
rect -120 780 -108 792
rect -96 780 -84 792
rect -72 780 -60 792
rect -48 780 -36 792
rect -24 780 -12 792
rect 0 780 12 792
rect 24 780 36 792
rect 48 780 60 792
rect 72 780 84 792
rect 96 780 108 792
rect 120 780 132 792
rect 144 780 156 792
rect 168 780 180 792
rect 192 780 204 792
rect 216 780 228 792
rect 240 780 252 792
rect 264 780 276 792
rect 288 780 300 792
rect 312 780 324 792
rect 336 780 348 792
rect 360 780 372 792
rect 384 780 396 792
rect 408 780 420 792
rect 432 780 444 792
rect 456 780 468 792
rect 480 780 492 792
rect 504 780 516 792
rect 528 780 540 792
rect 552 780 564 792
rect 576 780 588 792
rect 600 780 612 792
rect 624 780 636 792
rect 648 780 660 792
rect 672 780 684 792
rect 696 780 708 792
rect 720 780 732 792
rect 744 780 756 792
rect 768 780 780 792
rect 792 780 804 792
rect 816 780 828 792
rect 840 780 852 792
rect 864 780 876 792
rect 888 780 900 792
rect 912 780 924 792
rect 936 780 948 792
rect 960 780 972 792
rect 984 780 996 792
rect 1008 780 1020 792
rect 1032 780 1044 792
rect 1056 780 1068 792
rect 1080 780 1092 792
rect 1104 780 1116 792
rect 1128 780 1140 792
rect 1152 780 1164 792
rect 1176 780 1188 792
rect 1200 780 1212 792
rect 1224 780 1236 792
rect 1248 780 1260 792
rect 1272 780 1284 792
rect 1296 780 1308 792
rect 1320 780 1332 792
rect 1344 780 1356 792
rect 1368 780 1380 792
rect 1392 780 1404 792
rect 1416 780 1428 792
rect 1440 780 1452 792
rect 1464 780 1476 792
rect 1488 780 1500 792
rect 1512 780 1524 792
rect 1536 780 1548 792
rect 1560 780 1572 792
rect 1584 780 1596 792
rect 1608 780 1620 792
rect 1632 780 1644 792
rect 1656 780 1668 792
rect 1680 780 1692 792
rect 1704 780 1716 792
rect 1728 780 1740 792
rect 1752 780 1764 792
rect 1776 780 1788 792
rect 1800 780 1812 792
rect 1824 780 1836 792
rect 1848 780 1860 792
rect 1872 780 1884 792
rect 1896 780 1908 792
rect 1920 780 1932 792
rect 1944 780 1956 792
rect 1968 780 1980 792
rect 1992 780 2004 792
rect 2016 780 2028 792
rect 2040 780 2052 792
rect 2064 780 2076 792
rect 2088 780 2100 792
rect 2112 780 2124 792
rect 2136 780 2148 792
rect 2160 780 2172 792
rect 2184 780 2196 792
rect 2208 780 2220 792
rect 2232 780 2244 792
rect 2256 780 2268 792
rect 2280 780 2292 792
rect 2304 780 2316 792
rect 2328 780 2340 792
rect 2352 780 2364 792
rect 2376 780 2388 792
rect 2400 780 2412 792
rect 2424 780 2436 792
rect 2448 780 2460 792
rect 2472 780 2484 792
rect 2496 780 2508 792
rect 2520 780 2532 792
rect 2544 780 2556 792
rect 2568 780 2580 792
rect 2592 780 2604 792
rect 2616 780 2628 792
rect 2640 780 2652 792
rect 2664 780 2676 792
rect 2688 780 2700 792
rect 2712 780 2724 792
rect 2736 780 2748 792
rect 2760 780 2772 792
rect 2784 780 2796 792
rect 2808 780 2820 792
rect 2832 780 2844 792
rect 2856 780 2868 792
rect 2880 780 2892 792
rect 2904 780 2916 792
rect 2928 780 2940 792
rect 2952 780 2988 792
rect -1020 756 2988 780
rect -1020 744 -996 756
rect -984 744 -972 756
rect -960 744 -948 756
rect -936 744 -924 756
rect -912 744 -900 756
rect -888 744 -876 756
rect -864 744 -852 756
rect -840 744 -828 756
rect -816 744 -804 756
rect -792 744 -780 756
rect -768 744 -756 756
rect -744 744 -732 756
rect -720 744 -708 756
rect -696 744 -684 756
rect -672 744 -660 756
rect -648 744 -636 756
rect -624 744 -612 756
rect -600 744 -588 756
rect -576 744 -564 756
rect -552 744 -540 756
rect -528 744 -516 756
rect -504 744 -492 756
rect -480 744 -468 756
rect -456 744 -444 756
rect -432 744 -420 756
rect -408 744 -396 756
rect -384 744 -372 756
rect -360 744 -348 756
rect -336 744 -324 756
rect -312 744 -300 756
rect -288 744 -276 756
rect -264 744 -252 756
rect -240 744 -228 756
rect -216 744 -204 756
rect -192 744 -180 756
rect -168 744 -156 756
rect -144 744 -132 756
rect -120 744 -108 756
rect -96 744 -84 756
rect -72 744 -60 756
rect -48 744 -36 756
rect -24 744 -12 756
rect 0 744 12 756
rect 24 744 36 756
rect 48 744 60 756
rect 72 744 84 756
rect 96 744 108 756
rect 120 744 132 756
rect 144 744 156 756
rect 168 744 180 756
rect 192 744 204 756
rect 216 744 228 756
rect 240 744 252 756
rect 264 744 276 756
rect 288 744 300 756
rect 312 744 324 756
rect 336 744 348 756
rect 360 744 372 756
rect 384 744 396 756
rect 408 744 420 756
rect 432 744 444 756
rect 456 744 468 756
rect 480 744 492 756
rect 504 744 516 756
rect 528 744 540 756
rect 552 744 564 756
rect 576 744 588 756
rect 600 744 612 756
rect 624 744 636 756
rect 648 744 660 756
rect 672 744 684 756
rect 696 744 708 756
rect 720 744 732 756
rect 744 744 756 756
rect 768 744 780 756
rect 792 744 804 756
rect 816 744 828 756
rect 840 744 852 756
rect 864 744 876 756
rect 888 744 900 756
rect 912 744 924 756
rect 936 744 948 756
rect 960 744 972 756
rect 984 744 996 756
rect 1008 744 1020 756
rect 1032 744 1044 756
rect 1056 744 1068 756
rect 1080 744 1092 756
rect 1104 744 1116 756
rect 1128 744 1140 756
rect 1152 744 1164 756
rect 1176 744 1188 756
rect 1200 744 1212 756
rect 1224 744 1236 756
rect 1248 744 1260 756
rect 1272 744 1284 756
rect 1296 744 1308 756
rect 1320 744 1332 756
rect 1344 744 1356 756
rect 1368 744 1380 756
rect 1392 744 1404 756
rect 1416 744 1428 756
rect 1440 744 1452 756
rect 1464 744 1476 756
rect 1488 744 1500 756
rect 1512 744 1524 756
rect 1536 744 1548 756
rect 1560 744 1572 756
rect 1584 744 1596 756
rect 1608 744 1620 756
rect 1632 744 1644 756
rect 1656 744 1668 756
rect 1680 744 1692 756
rect 1704 744 1716 756
rect 1728 744 1740 756
rect 1752 744 1764 756
rect 1776 744 1788 756
rect 1800 744 1812 756
rect 1824 744 1836 756
rect 1848 744 1860 756
rect 1872 744 1884 756
rect 1896 744 1908 756
rect 1920 744 1932 756
rect 1944 744 1956 756
rect 1968 744 1980 756
rect 1992 744 2004 756
rect 2016 744 2028 756
rect 2040 744 2052 756
rect 2064 744 2076 756
rect 2088 744 2100 756
rect 2112 744 2124 756
rect 2136 744 2148 756
rect 2160 744 2172 756
rect 2184 744 2196 756
rect 2208 744 2220 756
rect 2232 744 2244 756
rect 2256 744 2268 756
rect 2280 744 2292 756
rect 2304 744 2316 756
rect 2328 744 2340 756
rect 2352 744 2364 756
rect 2376 744 2388 756
rect 2400 744 2412 756
rect 2424 744 2436 756
rect 2448 744 2460 756
rect 2472 744 2484 756
rect 2496 744 2508 756
rect 2520 744 2532 756
rect 2544 744 2556 756
rect 2568 744 2580 756
rect 2592 744 2604 756
rect 2616 744 2628 756
rect 2640 744 2652 756
rect 2664 744 2676 756
rect 2688 744 2700 756
rect 2712 744 2724 756
rect 2736 744 2748 756
rect 2760 744 2772 756
rect 2784 744 2796 756
rect 2808 744 2820 756
rect 2832 744 2844 756
rect 2856 744 2868 756
rect 2880 744 2892 756
rect 2904 744 2916 756
rect 2928 744 2940 756
rect 2952 744 2988 756
rect -1020 720 2988 744
rect -1020 708 -996 720
rect -984 708 -972 720
rect -960 708 -948 720
rect -936 708 -924 720
rect -912 708 -900 720
rect -888 708 -876 720
rect -864 708 -852 720
rect -840 708 -828 720
rect -816 708 -804 720
rect -792 708 -780 720
rect -768 708 -756 720
rect -744 708 -732 720
rect -720 708 -708 720
rect -696 708 -684 720
rect -672 708 -660 720
rect -648 708 -636 720
rect -624 708 -612 720
rect -600 708 -588 720
rect -576 708 -564 720
rect -552 708 -540 720
rect -528 708 -516 720
rect -504 708 -492 720
rect -480 708 -468 720
rect -456 708 -444 720
rect -432 708 -420 720
rect -408 708 -396 720
rect -384 708 -372 720
rect -360 708 -348 720
rect -336 708 -324 720
rect -312 708 -300 720
rect -288 708 -276 720
rect -264 708 -252 720
rect -240 708 -228 720
rect -216 708 -204 720
rect -192 708 -180 720
rect -168 708 -156 720
rect -144 708 -132 720
rect -120 708 -108 720
rect -96 708 -84 720
rect -72 708 -60 720
rect -48 708 -36 720
rect -24 708 -12 720
rect 0 708 12 720
rect 24 708 36 720
rect 48 708 60 720
rect 72 708 84 720
rect 96 708 108 720
rect 120 708 132 720
rect 144 708 156 720
rect 168 708 180 720
rect 192 708 204 720
rect 216 708 228 720
rect 240 708 252 720
rect 264 708 276 720
rect 288 708 300 720
rect 312 708 324 720
rect 336 708 348 720
rect 360 708 372 720
rect 384 708 396 720
rect 408 708 420 720
rect 432 708 444 720
rect 456 708 468 720
rect 480 708 492 720
rect 504 708 516 720
rect 528 708 540 720
rect 552 708 564 720
rect 576 708 588 720
rect 600 708 612 720
rect 624 708 636 720
rect 648 708 660 720
rect 672 708 684 720
rect 696 708 708 720
rect 720 708 732 720
rect 744 708 756 720
rect 768 708 780 720
rect 792 708 804 720
rect 816 708 828 720
rect 840 708 852 720
rect 864 708 876 720
rect 888 708 900 720
rect 912 708 924 720
rect 936 708 948 720
rect 960 708 972 720
rect 984 708 996 720
rect 1008 708 1020 720
rect 1032 708 1044 720
rect 1056 708 1068 720
rect 1080 708 1092 720
rect 1104 708 1116 720
rect 1128 708 1140 720
rect 1152 708 1164 720
rect 1176 708 1188 720
rect 1200 708 1212 720
rect 1224 708 1236 720
rect 1248 708 1260 720
rect 1272 708 1284 720
rect 1296 708 1308 720
rect 1320 708 1332 720
rect 1344 708 1356 720
rect 1368 708 1380 720
rect 1392 708 1404 720
rect 1416 708 1428 720
rect 1440 708 1452 720
rect 1464 708 1476 720
rect 1488 708 1500 720
rect 1512 708 1524 720
rect 1536 708 1548 720
rect 1560 708 1572 720
rect 1584 708 1596 720
rect 1608 708 1620 720
rect 1632 708 1644 720
rect 1656 708 1668 720
rect 1680 708 1692 720
rect 1704 708 1716 720
rect 1728 708 1740 720
rect 1752 708 1764 720
rect 1776 708 1788 720
rect 1800 708 1812 720
rect 1824 708 1836 720
rect 1848 708 1860 720
rect 1872 708 1884 720
rect 1896 708 1908 720
rect 1920 708 1932 720
rect 1944 708 1956 720
rect 1968 708 1980 720
rect 1992 708 2004 720
rect 2016 708 2028 720
rect 2040 708 2052 720
rect 2064 708 2076 720
rect 2088 708 2100 720
rect 2112 708 2124 720
rect 2136 708 2148 720
rect 2160 708 2172 720
rect 2184 708 2196 720
rect 2208 708 2220 720
rect 2232 708 2244 720
rect 2256 708 2268 720
rect 2280 708 2292 720
rect 2304 708 2316 720
rect 2328 708 2340 720
rect 2352 708 2364 720
rect 2376 708 2388 720
rect 2400 708 2412 720
rect 2424 708 2436 720
rect 2448 708 2460 720
rect 2472 708 2484 720
rect 2496 708 2508 720
rect 2520 708 2532 720
rect 2544 708 2556 720
rect 2568 708 2580 720
rect 2592 708 2604 720
rect 2616 708 2628 720
rect 2640 708 2652 720
rect 2664 708 2676 720
rect 2688 708 2700 720
rect 2712 708 2724 720
rect 2736 708 2748 720
rect 2760 708 2772 720
rect 2784 708 2796 720
rect 2808 708 2820 720
rect 2832 708 2844 720
rect 2856 708 2868 720
rect 2880 708 2892 720
rect 2904 708 2916 720
rect 2928 708 2940 720
rect 2952 708 2988 720
rect -1020 684 2988 708
rect -1020 672 -996 684
rect -984 672 -972 684
rect -960 672 -948 684
rect -936 672 -924 684
rect -912 672 -900 684
rect -888 672 -876 684
rect -864 672 -852 684
rect -840 672 -828 684
rect -816 672 -804 684
rect -792 672 -780 684
rect -768 672 -756 684
rect -744 672 -732 684
rect -720 672 -708 684
rect -696 672 -684 684
rect -672 672 -660 684
rect -648 672 -636 684
rect -624 672 -612 684
rect -600 672 -588 684
rect -576 672 -564 684
rect -552 672 -540 684
rect -528 672 -516 684
rect -504 672 -492 684
rect -480 672 -468 684
rect -456 672 -444 684
rect -432 672 -420 684
rect -408 672 -396 684
rect -384 672 -372 684
rect -360 672 -348 684
rect -336 672 -324 684
rect -312 672 -300 684
rect -288 672 -276 684
rect -264 672 -252 684
rect -240 672 -228 684
rect -216 672 -204 684
rect -192 672 -180 684
rect -168 672 -156 684
rect -144 672 -132 684
rect -120 672 -108 684
rect -96 672 -84 684
rect -72 672 -60 684
rect -48 672 -36 684
rect -24 672 -12 684
rect 0 672 12 684
rect 24 672 36 684
rect 48 672 60 684
rect 72 672 84 684
rect 96 672 108 684
rect 120 672 132 684
rect 144 672 156 684
rect 168 672 180 684
rect 192 672 204 684
rect 216 672 228 684
rect 240 672 252 684
rect 264 672 276 684
rect 288 672 300 684
rect 312 672 324 684
rect 336 672 348 684
rect 360 672 372 684
rect 384 672 396 684
rect 408 672 420 684
rect 432 672 444 684
rect 456 672 468 684
rect 480 672 492 684
rect 504 672 516 684
rect 528 672 540 684
rect 552 672 564 684
rect 576 672 588 684
rect 600 672 612 684
rect 624 672 636 684
rect 648 672 660 684
rect 672 672 684 684
rect 696 672 708 684
rect 720 672 732 684
rect 744 672 756 684
rect 768 672 780 684
rect 792 672 804 684
rect 816 672 828 684
rect 840 672 852 684
rect 864 672 876 684
rect 888 672 900 684
rect 912 672 924 684
rect 936 672 948 684
rect 960 672 972 684
rect 984 672 996 684
rect 1008 672 1020 684
rect 1032 672 1044 684
rect 1056 672 1068 684
rect 1080 672 1092 684
rect 1104 672 1116 684
rect 1128 672 1140 684
rect 1152 672 1164 684
rect 1176 672 1188 684
rect 1200 672 1212 684
rect 1224 672 1236 684
rect 1248 672 1260 684
rect 1272 672 1284 684
rect 1296 672 1308 684
rect 1320 672 1332 684
rect 1344 672 1356 684
rect 1368 672 1380 684
rect 1392 672 1404 684
rect 1416 672 1428 684
rect 1440 672 1452 684
rect 1464 672 1476 684
rect 1488 672 1500 684
rect 1512 672 1524 684
rect 1536 672 1548 684
rect 1560 672 1572 684
rect 1584 672 1596 684
rect 1608 672 1620 684
rect 1632 672 1644 684
rect 1656 672 1668 684
rect 1680 672 1692 684
rect 1704 672 1716 684
rect 1728 672 1740 684
rect 1752 672 1764 684
rect 1776 672 1788 684
rect 1800 672 1812 684
rect 1824 672 1836 684
rect 1848 672 1860 684
rect 1872 672 1884 684
rect 1896 672 1908 684
rect 1920 672 1932 684
rect 1944 672 1956 684
rect 1968 672 1980 684
rect 1992 672 2004 684
rect 2016 672 2028 684
rect 2040 672 2052 684
rect 2064 672 2076 684
rect 2088 672 2100 684
rect 2112 672 2124 684
rect 2136 672 2148 684
rect 2160 672 2172 684
rect 2184 672 2196 684
rect 2208 672 2220 684
rect 2232 672 2244 684
rect 2256 672 2268 684
rect 2280 672 2292 684
rect 2304 672 2316 684
rect 2328 672 2340 684
rect 2352 672 2364 684
rect 2376 672 2388 684
rect 2400 672 2412 684
rect 2424 672 2436 684
rect 2448 672 2460 684
rect 2472 672 2484 684
rect 2496 672 2508 684
rect 2520 672 2532 684
rect 2544 672 2556 684
rect 2568 672 2580 684
rect 2592 672 2604 684
rect 2616 672 2628 684
rect 2640 672 2652 684
rect 2664 672 2676 684
rect 2688 672 2700 684
rect 2712 672 2724 684
rect 2736 672 2748 684
rect 2760 672 2772 684
rect 2784 672 2796 684
rect 2808 672 2820 684
rect 2832 672 2844 684
rect 2856 672 2868 684
rect 2880 672 2892 684
rect 2904 672 2916 684
rect 2928 672 2940 684
rect 2952 672 2988 684
rect -1020 660 2988 672
rect -1116 648 -1104 660
rect -1092 648 -1056 660
rect -1044 648 2988 660
rect -1116 624 -1080 636
rect -1068 624 -1008 636
rect -996 624 -984 636
rect -972 624 -960 636
rect -948 624 -936 636
rect -924 624 -912 636
rect -900 624 -888 636
rect -876 624 -864 636
rect -852 624 -840 636
rect -828 624 -804 636
rect -792 624 -780 636
rect -768 624 -756 636
rect -744 624 -732 636
rect -720 624 -708 636
rect -696 624 -684 636
rect -672 624 -660 636
rect -648 624 -636 636
rect -624 624 -612 636
rect -600 624 -588 636
rect -576 624 -564 636
rect -552 624 -540 636
rect -528 624 -516 636
rect -504 624 -492 636
rect -480 624 -468 636
rect -456 624 -444 636
rect -432 624 -408 636
rect -396 624 -384 636
rect -372 624 -360 636
rect -348 624 -336 636
rect -324 624 -312 636
rect -300 624 -288 636
rect -276 624 -264 636
rect -252 624 -240 636
rect -228 624 -204 636
rect -192 624 -180 636
rect -168 624 -156 636
rect -144 624 -132 636
rect -120 624 -108 636
rect -96 624 -84 636
rect -72 624 -60 636
rect -48 624 -36 636
rect -24 624 -12 636
rect 0 624 12 636
rect 24 624 36 636
rect 48 624 60 636
rect 72 624 84 636
rect 96 624 108 636
rect 120 624 132 636
rect 144 624 156 636
rect 168 624 180 636
rect 192 624 204 636
rect 216 624 228 636
rect 240 624 252 636
rect 264 624 276 636
rect 288 624 300 636
rect 312 624 324 636
rect 336 624 348 636
rect 360 624 384 636
rect 396 624 408 636
rect 420 624 432 636
rect 444 624 456 636
rect 468 624 480 636
rect 492 624 504 636
rect 516 624 528 636
rect 540 624 552 636
rect 564 624 576 636
rect 588 624 600 636
rect 612 624 624 636
rect 636 624 648 636
rect 660 624 672 636
rect 684 624 696 636
rect 708 624 720 636
rect 732 624 744 636
rect 756 624 768 636
rect 780 624 792 636
rect 804 624 816 636
rect 828 624 840 636
rect 852 624 864 636
rect 876 624 888 636
rect 900 624 912 636
rect 924 624 936 636
rect 948 624 972 636
rect 984 624 996 636
rect 1008 624 1020 636
rect 1032 624 1044 636
rect 1056 624 1068 636
rect 1080 624 1092 636
rect 1104 624 1116 636
rect 1128 624 1140 636
rect 1152 624 1164 636
rect 1176 624 1188 636
rect 1200 624 1212 636
rect 1224 624 1236 636
rect 1248 624 1260 636
rect 1272 624 1284 636
rect 1296 624 1308 636
rect 1320 624 1332 636
rect 1344 624 1356 636
rect 1368 624 1380 636
rect 1392 624 1404 636
rect 1416 624 1428 636
rect 1440 624 1452 636
rect 1464 624 1476 636
rect 1488 624 1500 636
rect 1512 624 1524 636
rect 1536 624 1560 636
rect 1572 624 1584 636
rect 1596 624 1608 636
rect 1620 624 1632 636
rect 1644 624 1656 636
rect 1668 624 1680 636
rect 1692 624 1704 636
rect 1716 624 1728 636
rect 1740 624 1752 636
rect 1764 624 1776 636
rect 1788 624 1800 636
rect 1812 624 1824 636
rect 1836 624 1848 636
rect 1860 624 1872 636
rect 1884 624 1896 636
rect 1908 624 1920 636
rect 1932 624 1956 636
rect 1968 624 1980 636
rect 1992 624 2004 636
rect 2016 624 2028 636
rect 2040 624 2052 636
rect 2064 624 2076 636
rect 2088 624 2100 636
rect 2112 624 2124 636
rect 2136 624 2160 636
rect 2172 624 2184 636
rect 2196 624 2208 636
rect 2220 624 2232 636
rect 2244 624 2256 636
rect 2268 624 2280 636
rect 2292 624 2304 636
rect 2316 624 2328 636
rect 2340 624 2352 636
rect 2364 624 2376 636
rect 2388 624 2400 636
rect 2412 624 2424 636
rect 2436 624 2448 636
rect 2460 624 2472 636
rect 2484 624 2496 636
rect 2508 624 2520 636
rect 2532 624 2544 636
rect 2556 624 2568 636
rect 2580 624 2592 636
rect 2604 624 2616 636
rect 2628 624 2640 636
rect 2652 624 2664 636
rect 2676 624 2688 636
rect 2700 624 2712 636
rect 2724 624 2748 636
rect 2760 624 2772 636
rect 2784 624 2796 636
rect 2808 624 2820 636
rect 2832 624 2844 636
rect 2856 624 2868 636
rect 2880 624 2892 636
rect 2904 624 2916 636
rect 2928 624 2940 636
rect 2952 624 2964 636
rect 2976 624 2988 636
rect -1116 600 -1104 612
rect -1092 600 -1056 612
rect -1044 600 2988 612
rect -1116 -192 -1104 -180
rect -1092 -192 -1056 -180
rect -1044 -192 2988 -180
rect -1116 -216 -1080 -204
rect -1068 -216 -1008 -204
rect -996 -216 -984 -204
rect -972 -216 -960 -204
rect -948 -216 -936 -204
rect -924 -216 -912 -204
rect -900 -216 -888 -204
rect -876 -216 -864 -204
rect -852 -216 -840 -204
rect -828 -216 -804 -204
rect -792 -216 -780 -204
rect -768 -216 -756 -204
rect -744 -216 -732 -204
rect -720 -216 -708 -204
rect -696 -216 -684 -204
rect -672 -216 -660 -204
rect -648 -216 -636 -204
rect -624 -216 -612 -204
rect -600 -216 -588 -204
rect -576 -216 -564 -204
rect -552 -216 -540 -204
rect -528 -216 -516 -204
rect -504 -216 -492 -204
rect -480 -216 -468 -204
rect -456 -216 -444 -204
rect -432 -216 -408 -204
rect -396 -216 -384 -204
rect -372 -216 -360 -204
rect -348 -216 -336 -204
rect -324 -216 -312 -204
rect -300 -216 -288 -204
rect -276 -216 -264 -204
rect -252 -216 -240 -204
rect -228 -216 -204 -204
rect -192 -216 -180 -204
rect -168 -216 -156 -204
rect -144 -216 -132 -204
rect -120 -216 -108 -204
rect -96 -216 -84 -204
rect -72 -216 -60 -204
rect -48 -216 -36 -204
rect -24 -216 -12 -204
rect 0 -216 12 -204
rect 24 -216 36 -204
rect 48 -216 60 -204
rect 72 -216 84 -204
rect 96 -216 108 -204
rect 120 -216 132 -204
rect 144 -216 156 -204
rect 168 -216 180 -204
rect 192 -216 204 -204
rect 216 -216 228 -204
rect 240 -216 252 -204
rect 264 -216 276 -204
rect 288 -216 300 -204
rect 312 -216 324 -204
rect 336 -216 348 -204
rect 360 -216 384 -204
rect 396 -216 408 -204
rect 420 -216 432 -204
rect 444 -216 456 -204
rect 468 -216 480 -204
rect 492 -216 504 -204
rect 516 -216 528 -204
rect 540 -216 552 -204
rect 564 -216 576 -204
rect 588 -216 600 -204
rect 612 -216 624 -204
rect 636 -216 648 -204
rect 660 -216 672 -204
rect 684 -216 696 -204
rect 708 -216 720 -204
rect 732 -216 744 -204
rect 756 -216 768 -204
rect 780 -216 792 -204
rect 804 -216 816 -204
rect 828 -216 840 -204
rect 852 -216 864 -204
rect 876 -216 888 -204
rect 900 -216 912 -204
rect 924 -216 936 -204
rect 948 -216 972 -204
rect 984 -216 996 -204
rect 1008 -216 1020 -204
rect 1032 -216 1044 -204
rect 1056 -216 1068 -204
rect 1080 -216 1092 -204
rect 1104 -216 1116 -204
rect 1128 -216 1140 -204
rect 1152 -216 1164 -204
rect 1176 -216 1188 -204
rect 1200 -216 1212 -204
rect 1224 -216 1236 -204
rect 1248 -216 1260 -204
rect 1272 -216 1284 -204
rect 1296 -216 1308 -204
rect 1320 -216 1332 -204
rect 1344 -216 1356 -204
rect 1368 -216 1380 -204
rect 1392 -216 1404 -204
rect 1416 -216 1428 -204
rect 1440 -216 1452 -204
rect 1464 -216 1476 -204
rect 1488 -216 1500 -204
rect 1512 -216 1524 -204
rect 1536 -216 1560 -204
rect 1572 -216 1584 -204
rect 1596 -216 1608 -204
rect 1620 -216 1632 -204
rect 1644 -216 1656 -204
rect 1668 -216 1680 -204
rect 1692 -216 1704 -204
rect 1716 -216 1728 -204
rect 1740 -216 1752 -204
rect 1764 -216 1776 -204
rect 1788 -216 1800 -204
rect 1812 -216 1824 -204
rect 1836 -216 1848 -204
rect 1860 -216 1872 -204
rect 1884 -216 1896 -204
rect 1908 -216 1920 -204
rect 1932 -216 1956 -204
rect 1968 -216 1980 -204
rect 1992 -216 2004 -204
rect 2016 -216 2028 -204
rect 2040 -216 2052 -204
rect 2064 -216 2076 -204
rect 2088 -216 2100 -204
rect 2112 -216 2124 -204
rect 2136 -216 2160 -204
rect 2172 -216 2184 -204
rect 2196 -216 2208 -204
rect 2220 -216 2232 -204
rect 2244 -216 2256 -204
rect 2268 -216 2280 -204
rect 2292 -216 2304 -204
rect 2316 -216 2328 -204
rect 2340 -216 2352 -204
rect 2364 -216 2376 -204
rect 2388 -216 2400 -204
rect 2412 -216 2424 -204
rect 2436 -216 2448 -204
rect 2460 -216 2472 -204
rect 2484 -216 2496 -204
rect 2508 -216 2520 -204
rect 2532 -216 2544 -204
rect 2556 -216 2568 -204
rect 2580 -216 2592 -204
rect 2604 -216 2616 -204
rect 2628 -216 2640 -204
rect 2652 -216 2664 -204
rect 2676 -216 2688 -204
rect 2700 -216 2712 -204
rect 2724 -216 2748 -204
rect 2760 -216 2772 -204
rect 2784 -216 2796 -204
rect 2808 -216 2820 -204
rect 2832 -216 2844 -204
rect 2856 -216 2868 -204
rect 2880 -216 2892 -204
rect 2904 -216 2916 -204
rect 2928 -216 2940 -204
rect 2952 -216 2964 -204
rect 2976 -216 2988 -204
rect -1116 -240 -1104 -228
rect -1092 -240 -1056 -228
rect -1044 -240 2988 -228
rect -1020 -252 2988 -240
rect -1020 -264 -996 -252
rect -984 -264 -972 -252
rect -960 -264 -948 -252
rect -936 -264 -924 -252
rect -912 -264 -900 -252
rect -888 -264 -876 -252
rect -864 -264 -852 -252
rect -840 -264 -828 -252
rect -816 -264 -804 -252
rect -792 -264 -780 -252
rect -768 -264 -756 -252
rect -744 -264 -732 -252
rect -720 -264 -708 -252
rect -696 -264 -684 -252
rect -672 -264 -660 -252
rect -648 -264 -636 -252
rect -624 -264 -612 -252
rect -600 -264 -588 -252
rect -576 -264 -564 -252
rect -552 -264 -540 -252
rect -528 -264 -516 -252
rect -504 -264 -492 -252
rect -480 -264 -468 -252
rect -456 -264 -444 -252
rect -432 -264 -420 -252
rect -408 -264 -396 -252
rect -384 -264 -372 -252
rect -360 -264 -348 -252
rect -336 -264 -324 -252
rect -312 -264 -300 -252
rect -288 -264 -276 -252
rect -264 -264 -252 -252
rect -240 -264 -228 -252
rect -216 -264 -204 -252
rect -192 -264 -180 -252
rect -168 -264 -156 -252
rect -144 -264 -132 -252
rect -120 -264 -108 -252
rect -96 -264 -84 -252
rect -72 -264 -60 -252
rect -48 -264 -36 -252
rect -24 -264 -12 -252
rect 0 -264 12 -252
rect 24 -264 36 -252
rect 48 -264 60 -252
rect 72 -264 84 -252
rect 96 -264 108 -252
rect 120 -264 132 -252
rect 144 -264 156 -252
rect 168 -264 180 -252
rect 192 -264 204 -252
rect 216 -264 228 -252
rect 240 -264 252 -252
rect 264 -264 276 -252
rect 288 -264 300 -252
rect 312 -264 324 -252
rect 336 -264 348 -252
rect 360 -264 372 -252
rect 384 -264 396 -252
rect 408 -264 420 -252
rect 432 -264 444 -252
rect 456 -264 468 -252
rect 480 -264 492 -252
rect 504 -264 516 -252
rect 528 -264 540 -252
rect 552 -264 564 -252
rect 576 -264 588 -252
rect 600 -264 612 -252
rect 624 -264 636 -252
rect 648 -264 660 -252
rect 672 -264 684 -252
rect 696 -264 708 -252
rect 720 -264 732 -252
rect 744 -264 756 -252
rect 768 -264 780 -252
rect 792 -264 804 -252
rect 816 -264 828 -252
rect 840 -264 852 -252
rect 864 -264 876 -252
rect 888 -264 900 -252
rect 912 -264 924 -252
rect 936 -264 948 -252
rect 960 -264 972 -252
rect 984 -264 996 -252
rect 1008 -264 1020 -252
rect 1032 -264 1044 -252
rect 1056 -264 1068 -252
rect 1080 -264 1092 -252
rect 1104 -264 1116 -252
rect 1128 -264 1140 -252
rect 1152 -264 1164 -252
rect 1176 -264 1188 -252
rect 1200 -264 1212 -252
rect 1224 -264 1236 -252
rect 1248 -264 1260 -252
rect 1272 -264 1284 -252
rect 1296 -264 1308 -252
rect 1320 -264 1332 -252
rect 1344 -264 1356 -252
rect 1368 -264 1380 -252
rect 1392 -264 1404 -252
rect 1416 -264 1428 -252
rect 1440 -264 1452 -252
rect 1464 -264 1476 -252
rect 1488 -264 1500 -252
rect 1512 -264 1524 -252
rect 1536 -264 1548 -252
rect 1560 -264 1572 -252
rect 1584 -264 1596 -252
rect 1608 -264 1620 -252
rect 1632 -264 1644 -252
rect 1656 -264 1668 -252
rect 1680 -264 1692 -252
rect 1704 -264 1716 -252
rect 1728 -264 1740 -252
rect 1752 -264 1764 -252
rect 1776 -264 1788 -252
rect 1800 -264 1812 -252
rect 1824 -264 1836 -252
rect 1848 -264 1860 -252
rect 1872 -264 1884 -252
rect 1896 -264 1908 -252
rect 1920 -264 1932 -252
rect 1944 -264 1956 -252
rect 1968 -264 1980 -252
rect 1992 -264 2004 -252
rect 2016 -264 2028 -252
rect 2040 -264 2052 -252
rect 2064 -264 2076 -252
rect 2088 -264 2100 -252
rect 2112 -264 2124 -252
rect 2136 -264 2148 -252
rect 2160 -264 2172 -252
rect 2184 -264 2196 -252
rect 2208 -264 2220 -252
rect 2232 -264 2244 -252
rect 2256 -264 2268 -252
rect 2280 -264 2292 -252
rect 2304 -264 2316 -252
rect 2328 -264 2340 -252
rect 2352 -264 2364 -252
rect 2376 -264 2388 -252
rect 2400 -264 2412 -252
rect 2424 -264 2436 -252
rect 2448 -264 2460 -252
rect 2472 -264 2484 -252
rect 2496 -264 2508 -252
rect 2520 -264 2532 -252
rect 2544 -264 2556 -252
rect 2568 -264 2580 -252
rect 2592 -264 2604 -252
rect 2616 -264 2628 -252
rect 2640 -264 2652 -252
rect 2664 -264 2676 -252
rect 2688 -264 2700 -252
rect 2712 -264 2724 -252
rect 2736 -264 2748 -252
rect 2760 -264 2772 -252
rect 2784 -264 2796 -252
rect 2808 -264 2820 -252
rect 2832 -264 2844 -252
rect 2856 -264 2868 -252
rect 2880 -264 2892 -252
rect 2904 -264 2916 -252
rect 2928 -264 2940 -252
rect 2952 -264 2988 -252
rect -1020 -288 2988 -264
rect -1020 -300 -996 -288
rect -984 -300 -972 -288
rect -960 -300 -948 -288
rect -936 -300 -924 -288
rect -912 -300 -900 -288
rect -888 -300 -876 -288
rect -864 -300 -852 -288
rect -840 -300 -828 -288
rect -816 -300 -804 -288
rect -792 -300 -780 -288
rect -768 -300 -756 -288
rect -744 -300 -732 -288
rect -720 -300 -708 -288
rect -696 -300 -684 -288
rect -672 -300 -660 -288
rect -648 -300 -636 -288
rect -624 -300 -612 -288
rect -600 -300 -588 -288
rect -576 -300 -564 -288
rect -552 -300 -540 -288
rect -528 -300 -516 -288
rect -504 -300 -492 -288
rect -480 -300 -468 -288
rect -456 -300 -444 -288
rect -432 -300 -420 -288
rect -408 -300 -396 -288
rect -384 -300 -372 -288
rect -360 -300 -348 -288
rect -336 -300 -324 -288
rect -312 -300 -300 -288
rect -288 -300 -276 -288
rect -264 -300 -252 -288
rect -240 -300 -228 -288
rect -216 -300 -204 -288
rect -192 -300 -180 -288
rect -168 -300 -156 -288
rect -144 -300 -132 -288
rect -120 -300 -108 -288
rect -96 -300 -84 -288
rect -72 -300 -60 -288
rect -48 -300 -36 -288
rect -24 -300 -12 -288
rect 0 -300 12 -288
rect 24 -300 36 -288
rect 48 -300 60 -288
rect 72 -300 84 -288
rect 96 -300 108 -288
rect 120 -300 132 -288
rect 144 -300 156 -288
rect 168 -300 180 -288
rect 192 -300 204 -288
rect 216 -300 228 -288
rect 240 -300 252 -288
rect 264 -300 276 -288
rect 288 -300 300 -288
rect 312 -300 324 -288
rect 336 -300 348 -288
rect 360 -300 372 -288
rect 384 -300 396 -288
rect 408 -300 420 -288
rect 432 -300 444 -288
rect 456 -300 468 -288
rect 480 -300 492 -288
rect 504 -300 516 -288
rect 528 -300 540 -288
rect 552 -300 564 -288
rect 576 -300 588 -288
rect 600 -300 612 -288
rect 624 -300 636 -288
rect 648 -300 660 -288
rect 672 -300 684 -288
rect 696 -300 708 -288
rect 720 -300 732 -288
rect 744 -300 756 -288
rect 768 -300 780 -288
rect 792 -300 804 -288
rect 816 -300 828 -288
rect 840 -300 852 -288
rect 864 -300 876 -288
rect 888 -300 900 -288
rect 912 -300 924 -288
rect 936 -300 948 -288
rect 960 -300 972 -288
rect 984 -300 996 -288
rect 1008 -300 1020 -288
rect 1032 -300 1044 -288
rect 1056 -300 1068 -288
rect 1080 -300 1092 -288
rect 1104 -300 1116 -288
rect 1128 -300 1140 -288
rect 1152 -300 1164 -288
rect 1176 -300 1188 -288
rect 1200 -300 1212 -288
rect 1224 -300 1236 -288
rect 1248 -300 1260 -288
rect 1272 -300 1284 -288
rect 1296 -300 1308 -288
rect 1320 -300 1332 -288
rect 1344 -300 1356 -288
rect 1368 -300 1380 -288
rect 1392 -300 1404 -288
rect 1416 -300 1428 -288
rect 1440 -300 1452 -288
rect 1464 -300 1476 -288
rect 1488 -300 1500 -288
rect 1512 -300 1524 -288
rect 1536 -300 1548 -288
rect 1560 -300 1572 -288
rect 1584 -300 1596 -288
rect 1608 -300 1620 -288
rect 1632 -300 1644 -288
rect 1656 -300 1668 -288
rect 1680 -300 1692 -288
rect 1704 -300 1716 -288
rect 1728 -300 1740 -288
rect 1752 -300 1764 -288
rect 1776 -300 1788 -288
rect 1800 -300 1812 -288
rect 1824 -300 1836 -288
rect 1848 -300 1860 -288
rect 1872 -300 1884 -288
rect 1896 -300 1908 -288
rect 1920 -300 1932 -288
rect 1944 -300 1956 -288
rect 1968 -300 1980 -288
rect 1992 -300 2004 -288
rect 2016 -300 2028 -288
rect 2040 -300 2052 -288
rect 2064 -300 2076 -288
rect 2088 -300 2100 -288
rect 2112 -300 2124 -288
rect 2136 -300 2148 -288
rect 2160 -300 2172 -288
rect 2184 -300 2196 -288
rect 2208 -300 2220 -288
rect 2232 -300 2244 -288
rect 2256 -300 2268 -288
rect 2280 -300 2292 -288
rect 2304 -300 2316 -288
rect 2328 -300 2340 -288
rect 2352 -300 2364 -288
rect 2376 -300 2388 -288
rect 2400 -300 2412 -288
rect 2424 -300 2436 -288
rect 2448 -300 2460 -288
rect 2472 -300 2484 -288
rect 2496 -300 2508 -288
rect 2520 -300 2532 -288
rect 2544 -300 2556 -288
rect 2568 -300 2580 -288
rect 2592 -300 2604 -288
rect 2616 -300 2628 -288
rect 2640 -300 2652 -288
rect 2664 -300 2676 -288
rect 2688 -300 2700 -288
rect 2712 -300 2724 -288
rect 2736 -300 2748 -288
rect 2760 -300 2772 -288
rect 2784 -300 2796 -288
rect 2808 -300 2820 -288
rect 2832 -300 2844 -288
rect 2856 -300 2868 -288
rect 2880 -300 2892 -288
rect 2904 -300 2916 -288
rect 2928 -300 2940 -288
rect 2952 -300 2988 -288
rect -1020 -324 2988 -300
rect -1020 -336 -996 -324
rect -984 -336 -972 -324
rect -960 -336 -948 -324
rect -936 -336 -924 -324
rect -912 -336 -900 -324
rect -888 -336 -876 -324
rect -864 -336 -852 -324
rect -840 -336 -828 -324
rect -816 -336 -804 -324
rect -792 -336 -780 -324
rect -768 -336 -756 -324
rect -744 -336 -732 -324
rect -720 -336 -708 -324
rect -696 -336 -684 -324
rect -672 -336 -660 -324
rect -648 -336 -636 -324
rect -624 -336 -612 -324
rect -600 -336 -588 -324
rect -576 -336 -564 -324
rect -552 -336 -540 -324
rect -528 -336 -516 -324
rect -504 -336 -492 -324
rect -480 -336 -468 -324
rect -456 -336 -444 -324
rect -432 -336 -420 -324
rect -408 -336 -396 -324
rect -384 -336 -372 -324
rect -360 -336 -348 -324
rect -336 -336 -324 -324
rect -312 -336 -300 -324
rect -288 -336 -276 -324
rect -264 -336 -252 -324
rect -240 -336 -228 -324
rect -216 -336 -204 -324
rect -192 -336 -180 -324
rect -168 -336 -156 -324
rect -144 -336 -132 -324
rect -120 -336 -108 -324
rect -96 -336 -84 -324
rect -72 -336 -60 -324
rect -48 -336 -36 -324
rect -24 -336 -12 -324
rect 0 -336 12 -324
rect 24 -336 36 -324
rect 48 -336 60 -324
rect 72 -336 84 -324
rect 96 -336 108 -324
rect 120 -336 132 -324
rect 144 -336 156 -324
rect 168 -336 180 -324
rect 192 -336 204 -324
rect 216 -336 228 -324
rect 240 -336 252 -324
rect 264 -336 276 -324
rect 288 -336 300 -324
rect 312 -336 324 -324
rect 336 -336 348 -324
rect 360 -336 372 -324
rect 384 -336 396 -324
rect 408 -336 420 -324
rect 432 -336 444 -324
rect 456 -336 468 -324
rect 480 -336 492 -324
rect 504 -336 516 -324
rect 528 -336 540 -324
rect 552 -336 564 -324
rect 576 -336 588 -324
rect 600 -336 612 -324
rect 624 -336 636 -324
rect 648 -336 660 -324
rect 672 -336 684 -324
rect 696 -336 708 -324
rect 720 -336 732 -324
rect 744 -336 756 -324
rect 768 -336 780 -324
rect 792 -336 804 -324
rect 816 -336 828 -324
rect 840 -336 852 -324
rect 864 -336 876 -324
rect 888 -336 900 -324
rect 912 -336 924 -324
rect 936 -336 948 -324
rect 960 -336 972 -324
rect 984 -336 996 -324
rect 1008 -336 1020 -324
rect 1032 -336 1044 -324
rect 1056 -336 1068 -324
rect 1080 -336 1092 -324
rect 1104 -336 1116 -324
rect 1128 -336 1140 -324
rect 1152 -336 1164 -324
rect 1176 -336 1188 -324
rect 1200 -336 1212 -324
rect 1224 -336 1236 -324
rect 1248 -336 1260 -324
rect 1272 -336 1284 -324
rect 1296 -336 1308 -324
rect 1320 -336 1332 -324
rect 1344 -336 1356 -324
rect 1368 -336 1380 -324
rect 1392 -336 1404 -324
rect 1416 -336 1428 -324
rect 1440 -336 1452 -324
rect 1464 -336 1476 -324
rect 1488 -336 1500 -324
rect 1512 -336 1524 -324
rect 1536 -336 1548 -324
rect 1560 -336 1572 -324
rect 1584 -336 1596 -324
rect 1608 -336 1620 -324
rect 1632 -336 1644 -324
rect 1656 -336 1668 -324
rect 1680 -336 1692 -324
rect 1704 -336 1716 -324
rect 1728 -336 1740 -324
rect 1752 -336 1764 -324
rect 1776 -336 1788 -324
rect 1800 -336 1812 -324
rect 1824 -336 1836 -324
rect 1848 -336 1860 -324
rect 1872 -336 1884 -324
rect 1896 -336 1908 -324
rect 1920 -336 1932 -324
rect 1944 -336 1956 -324
rect 1968 -336 1980 -324
rect 1992 -336 2004 -324
rect 2016 -336 2028 -324
rect 2040 -336 2052 -324
rect 2064 -336 2076 -324
rect 2088 -336 2100 -324
rect 2112 -336 2124 -324
rect 2136 -336 2148 -324
rect 2160 -336 2172 -324
rect 2184 -336 2196 -324
rect 2208 -336 2220 -324
rect 2232 -336 2244 -324
rect 2256 -336 2268 -324
rect 2280 -336 2292 -324
rect 2304 -336 2316 -324
rect 2328 -336 2340 -324
rect 2352 -336 2364 -324
rect 2376 -336 2388 -324
rect 2400 -336 2412 -324
rect 2424 -336 2436 -324
rect 2448 -336 2460 -324
rect 2472 -336 2484 -324
rect 2496 -336 2508 -324
rect 2520 -336 2532 -324
rect 2544 -336 2556 -324
rect 2568 -336 2580 -324
rect 2592 -336 2604 -324
rect 2616 -336 2628 -324
rect 2640 -336 2652 -324
rect 2664 -336 2676 -324
rect 2688 -336 2700 -324
rect 2712 -336 2724 -324
rect 2736 -336 2748 -324
rect 2760 -336 2772 -324
rect 2784 -336 2796 -324
rect 2808 -336 2820 -324
rect 2832 -336 2844 -324
rect 2856 -336 2868 -324
rect 2880 -336 2892 -324
rect 2904 -336 2916 -324
rect 2928 -336 2940 -324
rect 2952 -336 2988 -324
rect -1020 -360 2988 -336
rect -1020 -372 -996 -360
rect -984 -372 -972 -360
rect -960 -372 -948 -360
rect -936 -372 -924 -360
rect -912 -372 -900 -360
rect -888 -372 -876 -360
rect -864 -372 -852 -360
rect -840 -372 -828 -360
rect -816 -372 -804 -360
rect -792 -372 -780 -360
rect -768 -372 -756 -360
rect -744 -372 -732 -360
rect -720 -372 -708 -360
rect -696 -372 -684 -360
rect -672 -372 -660 -360
rect -648 -372 -636 -360
rect -624 -372 -612 -360
rect -600 -372 -588 -360
rect -576 -372 -564 -360
rect -552 -372 -540 -360
rect -528 -372 -516 -360
rect -504 -372 -492 -360
rect -480 -372 -468 -360
rect -456 -372 -444 -360
rect -432 -372 -420 -360
rect -408 -372 -396 -360
rect -384 -372 -372 -360
rect -360 -372 -348 -360
rect -336 -372 -324 -360
rect -312 -372 -300 -360
rect -288 -372 -276 -360
rect -264 -372 -252 -360
rect -240 -372 -228 -360
rect -216 -372 -204 -360
rect -192 -372 -180 -360
rect -168 -372 -156 -360
rect -144 -372 -132 -360
rect -120 -372 -108 -360
rect -96 -372 -84 -360
rect -72 -372 -60 -360
rect -48 -372 -36 -360
rect -24 -372 -12 -360
rect 0 -372 12 -360
rect 24 -372 36 -360
rect 48 -372 60 -360
rect 72 -372 84 -360
rect 96 -372 108 -360
rect 120 -372 132 -360
rect 144 -372 156 -360
rect 168 -372 180 -360
rect 192 -372 204 -360
rect 216 -372 228 -360
rect 240 -372 252 -360
rect 264 -372 276 -360
rect 288 -372 300 -360
rect 312 -372 324 -360
rect 336 -372 348 -360
rect 360 -372 372 -360
rect 384 -372 396 -360
rect 408 -372 420 -360
rect 432 -372 444 -360
rect 456 -372 468 -360
rect 480 -372 492 -360
rect 504 -372 516 -360
rect 528 -372 540 -360
rect 552 -372 564 -360
rect 576 -372 588 -360
rect 600 -372 612 -360
rect 624 -372 636 -360
rect 648 -372 660 -360
rect 672 -372 684 -360
rect 696 -372 708 -360
rect 720 -372 732 -360
rect 744 -372 756 -360
rect 768 -372 780 -360
rect 792 -372 804 -360
rect 816 -372 828 -360
rect 840 -372 852 -360
rect 864 -372 876 -360
rect 888 -372 900 -360
rect 912 -372 924 -360
rect 936 -372 948 -360
rect 960 -372 972 -360
rect 984 -372 996 -360
rect 1008 -372 1020 -360
rect 1032 -372 1044 -360
rect 1056 -372 1068 -360
rect 1080 -372 1092 -360
rect 1104 -372 1116 -360
rect 1128 -372 1140 -360
rect 1152 -372 1164 -360
rect 1176 -372 1188 -360
rect 1200 -372 1212 -360
rect 1224 -372 1236 -360
rect 1248 -372 1260 -360
rect 1272 -372 1284 -360
rect 1296 -372 1308 -360
rect 1320 -372 1332 -360
rect 1344 -372 1356 -360
rect 1368 -372 1380 -360
rect 1392 -372 1404 -360
rect 1416 -372 1428 -360
rect 1440 -372 1452 -360
rect 1464 -372 1476 -360
rect 1488 -372 1500 -360
rect 1512 -372 1524 -360
rect 1536 -372 1548 -360
rect 1560 -372 1572 -360
rect 1584 -372 1596 -360
rect 1608 -372 1620 -360
rect 1632 -372 1644 -360
rect 1656 -372 1668 -360
rect 1680 -372 1692 -360
rect 1704 -372 1716 -360
rect 1728 -372 1740 -360
rect 1752 -372 1764 -360
rect 1776 -372 1788 -360
rect 1800 -372 1812 -360
rect 1824 -372 1836 -360
rect 1848 -372 1860 -360
rect 1872 -372 1884 -360
rect 1896 -372 1908 -360
rect 1920 -372 1932 -360
rect 1944 -372 1956 -360
rect 1968 -372 1980 -360
rect 1992 -372 2004 -360
rect 2016 -372 2028 -360
rect 2040 -372 2052 -360
rect 2064 -372 2076 -360
rect 2088 -372 2100 -360
rect 2112 -372 2124 -360
rect 2136 -372 2148 -360
rect 2160 -372 2172 -360
rect 2184 -372 2196 -360
rect 2208 -372 2220 -360
rect 2232 -372 2244 -360
rect 2256 -372 2268 -360
rect 2280 -372 2292 -360
rect 2304 -372 2316 -360
rect 2328 -372 2340 -360
rect 2352 -372 2364 -360
rect 2376 -372 2388 -360
rect 2400 -372 2412 -360
rect 2424 -372 2436 -360
rect 2448 -372 2460 -360
rect 2472 -372 2484 -360
rect 2496 -372 2508 -360
rect 2520 -372 2532 -360
rect 2544 -372 2556 -360
rect 2568 -372 2580 -360
rect 2592 -372 2604 -360
rect 2616 -372 2628 -360
rect 2640 -372 2652 -360
rect 2664 -372 2676 -360
rect 2688 -372 2700 -360
rect 2712 -372 2724 -360
rect 2736 -372 2748 -360
rect 2760 -372 2772 -360
rect 2784 -372 2796 -360
rect 2808 -372 2820 -360
rect 2832 -372 2844 -360
rect 2856 -372 2868 -360
rect 2880 -372 2892 -360
rect 2904 -372 2916 -360
rect 2928 -372 2940 -360
rect 2952 -372 2988 -360
rect -1020 -396 2988 -372
use nautanauta_cell  nautanauta_cell_0
timestamp 1665298770
transform 1 0 -228 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_1
timestamp 1665298770
transform 1 0 -108 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_2
timestamp 1665298770
transform 1 0 12 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_3
timestamp 1665298770
transform 1 0 132 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_4
timestamp 1665298770
transform 1 0 252 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_5
timestamp 1665298770
transform 1 0 372 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_6
timestamp 1665298770
transform 1 0 492 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_7
timestamp 1665298770
transform 1 0 612 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_8
timestamp 1665298770
transform 1 0 732 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_9
timestamp 1665298770
transform 1 0 852 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_10
timestamp 1665298770
transform -1 0 264 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_11
timestamp 1665298770
transform -1 0 144 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_12
timestamp 1665298770
transform -1 0 24 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_13
timestamp 1665298770
transform -1 0 -96 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_14
timestamp 1665298770
transform -1 0 -216 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_15
timestamp 1665298770
transform -1 0 -336 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_16
timestamp 1665298770
transform -1 0 2184 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_17
timestamp 1665298770
transform -1 0 2064 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_18
timestamp 1665298770
transform -1 0 1944 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_19
timestamp 1665298770
transform -1 0 1824 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_20
timestamp 1665298770
transform -1 0 1704 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_21
timestamp 1665298770
transform -1 0 1584 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_22
timestamp 1665298770
transform -1 0 1464 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_23
timestamp 1665298770
transform -1 0 1344 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_24
timestamp 1665298770
transform -1 0 1224 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_25
timestamp 1665298770
transform -1 0 1104 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_26
timestamp 1665298770
transform 1 0 2292 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_27
timestamp 1665298770
transform 1 0 2172 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_28
timestamp 1665298770
transform 1 0 2052 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_29
timestamp 1665298770
transform 1 0 1932 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_30
timestamp 1665298770
transform 1 0 1812 0 1 -36
box -720 -132 -588 612
use nautanauta_cell  nautanauta_cell_31
timestamp 1665298770
transform 1 0 1692 0 1 -36
box -720 -132 -588 612
use nautanauta_edge  nautanauta_edge_0
timestamp 1665298770
transform 1 0 -276 0 1 -36
box -756 -132 -660 612
use nautanauta_edge  nautanauta_edge_1
timestamp 1665298770
transform -1 0 2232 0 1 -36
box -756 -132 -660 612
<< labels >>
rlabel metal3 -1044 -168 -1032 -108 0 gnd
port 9 nsew
rlabel metal3 -1044 72 -1032 84 0 ip
port 1 nsew
rlabel metal3 -1044 120 -1032 132 0 im
port 2 nsew
rlabel metal3 -1044 240 -1032 252 0 op
port 3 nsew
rlabel metal3 -1044 -48 -1032 -36 0 om
port 4 nsew
rlabel metal3 -1044 492 -1032 552 0 vdd
port 5 nsew
rlabel metal3 -1044 420 -1032 432 0 gp
port 6 nsew
rlabel metal3 -1044 288 -1032 300 0 bp
port 7 nsew
rlabel metal3 -1044 444 -1032 456 0 vreg
port 8 nsew
rlabel metal3 -1044 204 -1032 216 0 xm
rlabel metal3 -1044 -12 -1032 0 0 xp
<< end >>
