magic
tech gf180mcuC
timestamp 1662387721
<< nwell >>
rect -48 246 180 372
rect -48 102 180 222
<< nmos >>
rect -24 -108 -12 -72
rect 0 -108 12 -72
rect 24 -108 36 -72
rect 48 -108 60 -72
rect 72 -108 84 -72
rect 96 -108 108 -72
rect 120 -108 132 -72
rect 144 -108 156 -72
<< pmos >>
rect -24 156 -12 186
rect 0 156 12 186
rect 24 156 36 186
rect 48 156 60 186
rect 72 156 84 186
rect 96 156 108 186
rect 120 156 132 186
rect 144 156 156 186
<< mvpmos >>
rect -24 300 -12 336
rect 0 300 12 336
rect 24 300 36 336
rect 48 300 60 336
rect 72 300 84 336
rect 96 300 108 336
rect 120 300 132 336
rect 144 300 156 336
<< ndiff >>
rect -36 -75 -24 -72
rect -36 -81 -33 -75
rect -27 -81 -24 -75
rect -36 -87 -24 -81
rect -36 -93 -33 -87
rect -27 -93 -24 -87
rect -36 -99 -24 -93
rect -36 -105 -33 -99
rect -27 -105 -24 -99
rect -36 -108 -24 -105
rect -12 -75 0 -72
rect -12 -81 -9 -75
rect -3 -81 0 -75
rect -12 -87 0 -81
rect -12 -93 -9 -87
rect -3 -93 0 -87
rect -12 -99 0 -93
rect -12 -105 -9 -99
rect -3 -105 0 -99
rect -12 -108 0 -105
rect 12 -75 24 -72
rect 12 -81 15 -75
rect 21 -81 24 -75
rect 12 -87 24 -81
rect 12 -93 15 -87
rect 21 -93 24 -87
rect 12 -99 24 -93
rect 12 -105 15 -99
rect 21 -105 24 -99
rect 12 -108 24 -105
rect 36 -75 48 -72
rect 36 -81 39 -75
rect 45 -81 48 -75
rect 36 -87 48 -81
rect 36 -93 39 -87
rect 45 -93 48 -87
rect 36 -99 48 -93
rect 36 -105 39 -99
rect 45 -105 48 -99
rect 36 -108 48 -105
rect 60 -75 72 -72
rect 60 -81 63 -75
rect 69 -81 72 -75
rect 60 -87 72 -81
rect 60 -93 63 -87
rect 69 -93 72 -87
rect 60 -99 72 -93
rect 60 -105 63 -99
rect 69 -105 72 -99
rect 60 -108 72 -105
rect 84 -75 96 -72
rect 84 -81 87 -75
rect 93 -81 96 -75
rect 84 -87 96 -81
rect 84 -93 87 -87
rect 93 -93 96 -87
rect 84 -99 96 -93
rect 84 -105 87 -99
rect 93 -105 96 -99
rect 84 -108 96 -105
rect 108 -75 120 -72
rect 108 -81 111 -75
rect 117 -81 120 -75
rect 108 -87 120 -81
rect 108 -93 111 -87
rect 117 -93 120 -87
rect 108 -99 120 -93
rect 108 -105 111 -99
rect 117 -105 120 -99
rect 108 -108 120 -105
rect 132 -75 144 -72
rect 132 -81 135 -75
rect 141 -81 144 -75
rect 132 -87 144 -81
rect 132 -93 135 -87
rect 141 -93 144 -87
rect 132 -99 144 -93
rect 132 -105 135 -99
rect 141 -105 144 -99
rect 132 -108 144 -105
rect 156 -75 168 -72
rect 156 -81 159 -75
rect 165 -81 168 -75
rect 156 -87 168 -81
rect 156 -93 159 -87
rect 165 -93 168 -87
rect 156 -99 168 -93
rect 156 -105 159 -99
rect 165 -105 168 -99
rect 156 -108 168 -105
<< pdiff >>
rect -36 177 -24 186
rect -36 171 -33 177
rect -27 171 -24 177
rect -36 165 -24 171
rect -36 159 -33 165
rect -27 159 -24 165
rect -36 156 -24 159
rect -12 177 0 186
rect -12 171 -9 177
rect -3 171 0 177
rect -12 165 0 171
rect -12 159 -9 165
rect -3 159 0 165
rect -12 156 0 159
rect 12 177 24 186
rect 12 171 15 177
rect 21 171 24 177
rect 12 165 24 171
rect 12 159 15 165
rect 21 159 24 165
rect 12 156 24 159
rect 36 177 48 186
rect 36 171 39 177
rect 45 171 48 177
rect 36 165 48 171
rect 36 159 39 165
rect 45 159 48 165
rect 36 156 48 159
rect 60 177 72 186
rect 60 171 63 177
rect 69 171 72 177
rect 60 165 72 171
rect 60 159 63 165
rect 69 159 72 165
rect 60 156 72 159
rect 84 177 96 186
rect 84 171 87 177
rect 93 171 96 177
rect 84 165 96 171
rect 84 159 87 165
rect 93 159 96 165
rect 84 156 96 159
rect 108 177 120 186
rect 108 171 111 177
rect 117 171 120 177
rect 108 165 120 171
rect 108 159 111 165
rect 117 159 120 165
rect 108 156 120 159
rect 132 177 144 186
rect 132 171 135 177
rect 141 171 144 177
rect 132 165 144 171
rect 132 159 135 165
rect 141 159 144 165
rect 132 156 144 159
rect 156 177 168 186
rect 156 171 159 177
rect 165 171 168 177
rect 156 165 168 171
rect 156 159 159 165
rect 165 159 168 165
rect 156 156 168 159
<< mvpdiff >>
rect -36 333 -24 336
rect -36 327 -33 333
rect -27 327 -24 333
rect -36 321 -24 327
rect -36 315 -33 321
rect -27 315 -24 321
rect -36 309 -24 315
rect -36 303 -33 309
rect -27 303 -24 309
rect -36 300 -24 303
rect -12 333 0 336
rect -12 327 -9 333
rect -3 327 0 333
rect -12 321 0 327
rect -12 315 -9 321
rect -3 315 0 321
rect -12 309 0 315
rect -12 303 -9 309
rect -3 303 0 309
rect -12 300 0 303
rect 12 333 24 336
rect 12 327 15 333
rect 21 327 24 333
rect 12 321 24 327
rect 12 315 15 321
rect 21 315 24 321
rect 12 309 24 315
rect 12 303 15 309
rect 21 303 24 309
rect 12 300 24 303
rect 36 333 48 336
rect 36 327 39 333
rect 45 327 48 333
rect 36 321 48 327
rect 36 315 39 321
rect 45 315 48 321
rect 36 309 48 315
rect 36 303 39 309
rect 45 303 48 309
rect 36 300 48 303
rect 60 333 72 336
rect 60 327 63 333
rect 69 327 72 333
rect 60 321 72 327
rect 60 315 63 321
rect 69 315 72 321
rect 60 309 72 315
rect 60 303 63 309
rect 69 303 72 309
rect 60 300 72 303
rect 84 333 96 336
rect 84 327 87 333
rect 93 327 96 333
rect 84 321 96 327
rect 84 315 87 321
rect 93 315 96 321
rect 84 309 96 315
rect 84 303 87 309
rect 93 303 96 309
rect 84 300 96 303
rect 108 333 120 336
rect 108 327 111 333
rect 117 327 120 333
rect 108 321 120 327
rect 108 315 111 321
rect 117 315 120 321
rect 108 309 120 315
rect 108 303 111 309
rect 117 303 120 309
rect 108 300 120 303
rect 132 333 144 336
rect 132 327 135 333
rect 141 327 144 333
rect 132 321 144 327
rect 132 315 135 321
rect 141 315 144 321
rect 132 309 144 315
rect 132 303 135 309
rect 141 303 144 309
rect 132 300 144 303
rect 156 333 168 336
rect 156 327 159 333
rect 165 327 168 333
rect 156 321 168 327
rect 156 315 159 321
rect 165 315 168 321
rect 156 309 168 315
rect 156 303 159 309
rect 165 303 168 309
rect 156 300 168 303
<< ndiffc >>
rect -33 -81 -27 -75
rect -33 -93 -27 -87
rect -33 -105 -27 -99
rect -9 -81 -3 -75
rect -9 -93 -3 -87
rect -9 -105 -3 -99
rect 15 -81 21 -75
rect 15 -93 21 -87
rect 15 -105 21 -99
rect 39 -81 45 -75
rect 39 -93 45 -87
rect 39 -105 45 -99
rect 63 -81 69 -75
rect 63 -93 69 -87
rect 63 -105 69 -99
rect 87 -81 93 -75
rect 87 -93 93 -87
rect 87 -105 93 -99
rect 111 -81 117 -75
rect 111 -93 117 -87
rect 111 -105 117 -99
rect 135 -81 141 -75
rect 135 -93 141 -87
rect 135 -105 141 -99
rect 159 -81 165 -75
rect 159 -93 165 -87
rect 159 -105 165 -99
<< pdiffc >>
rect -33 171 -27 177
rect -33 159 -27 165
rect -9 171 -3 177
rect -9 159 -3 165
rect 15 171 21 177
rect 15 159 21 165
rect 39 171 45 177
rect 39 159 45 165
rect 63 171 69 177
rect 63 159 69 165
rect 87 171 93 177
rect 87 159 93 165
rect 111 171 117 177
rect 111 159 117 165
rect 135 171 141 177
rect 135 159 141 165
rect 159 171 165 177
rect 159 159 165 165
<< mvpdiffc >>
rect -33 327 -27 333
rect -33 315 -27 321
rect -33 303 -27 309
rect -9 327 -3 333
rect -9 315 -3 321
rect -9 303 -3 309
rect 15 327 21 333
rect 15 315 21 321
rect 15 303 21 309
rect 39 327 45 333
rect 39 315 45 321
rect 39 303 45 309
rect 63 327 69 333
rect 63 315 69 321
rect 63 303 69 309
rect 87 327 93 333
rect 87 315 93 321
rect 87 303 93 309
rect 111 327 117 333
rect 111 315 117 321
rect 111 303 117 309
rect 135 327 141 333
rect 135 315 141 321
rect 135 303 141 309
rect 159 327 165 333
rect 159 315 165 321
rect 159 303 165 309
<< psubdiff >>
rect -48 405 180 408
rect -48 399 -45 405
rect -39 399 -33 405
rect -27 399 -21 405
rect -15 399 -9 405
rect -3 399 3 405
rect 9 399 15 405
rect 21 399 27 405
rect 33 399 39 405
rect 45 399 51 405
rect 57 399 63 405
rect 69 399 75 405
rect 81 399 87 405
rect 93 399 99 405
rect 105 399 111 405
rect 117 399 123 405
rect 129 399 135 405
rect 141 399 147 405
rect 153 399 159 405
rect 165 399 171 405
rect 177 399 180 405
rect -48 396 180 399
rect -48 237 180 240
rect -48 231 -45 237
rect -39 231 -33 237
rect -27 231 -21 237
rect -15 231 -9 237
rect -3 231 3 237
rect 9 231 15 237
rect 21 231 27 237
rect 33 231 39 237
rect 45 231 51 237
rect 57 231 63 237
rect 69 231 75 237
rect 81 231 87 237
rect 93 231 99 237
rect 105 231 111 237
rect 117 231 123 237
rect 129 231 135 237
rect 141 231 147 237
rect 153 231 159 237
rect 165 231 171 237
rect 177 231 180 237
rect -48 228 180 231
rect -48 45 180 48
rect -48 39 -45 45
rect -39 39 -33 45
rect -27 39 -21 45
rect -15 39 -9 45
rect -3 39 3 45
rect 9 39 15 45
rect 21 39 27 45
rect 33 39 39 45
rect 45 39 51 45
rect 57 39 63 45
rect 69 39 75 45
rect 81 39 87 45
rect 93 39 99 45
rect 105 39 111 45
rect 117 39 123 45
rect 129 39 135 45
rect 141 39 147 45
rect 153 39 159 45
rect 165 39 171 45
rect 177 39 180 45
rect -48 36 180 39
rect -48 -27 180 -24
rect -48 -33 -45 -27
rect -39 -33 -33 -27
rect -27 -33 -21 -27
rect -15 -33 -9 -27
rect -3 -33 3 -27
rect 9 -33 15 -27
rect 21 -33 27 -27
rect 33 -33 39 -27
rect 45 -33 51 -27
rect 57 -33 63 -27
rect 69 -33 75 -27
rect 81 -33 87 -27
rect 93 -33 99 -27
rect 105 -33 111 -27
rect 117 -33 123 -27
rect 129 -33 135 -27
rect 141 -33 147 -27
rect 153 -33 159 -27
rect 165 -33 171 -27
rect 177 -33 180 -27
rect -48 -36 180 -33
rect -48 -123 180 -120
rect -48 -129 -45 -123
rect -39 -129 -33 -123
rect -27 -129 -21 -123
rect -15 -129 -9 -123
rect -3 -129 3 -123
rect 9 -129 15 -123
rect 21 -129 27 -123
rect 33 -129 39 -123
rect 45 -129 51 -123
rect 57 -129 63 -123
rect 69 -129 75 -123
rect 81 -129 87 -123
rect 93 -129 99 -123
rect 105 -129 111 -123
rect 117 -129 123 -123
rect 129 -129 135 -123
rect 141 -129 147 -123
rect 153 -129 159 -123
rect 165 -129 171 -123
rect 177 -129 180 -123
rect -48 -132 180 -129
<< nsubdiff >>
rect -36 213 168 216
rect -36 207 -33 213
rect -27 207 -21 213
rect -15 207 -9 213
rect -3 207 3 213
rect 9 207 15 213
rect 21 207 27 213
rect 33 207 39 213
rect 45 207 51 213
rect 57 207 63 213
rect 69 207 75 213
rect 81 207 87 213
rect 93 207 99 213
rect 105 207 111 213
rect 117 207 123 213
rect 129 207 135 213
rect 141 207 147 213
rect 153 207 159 213
rect 165 207 168 213
rect -36 204 168 207
rect -36 117 168 120
rect -36 111 -33 117
rect -27 111 -21 117
rect -15 111 -9 117
rect -3 111 3 117
rect 9 111 15 117
rect 21 111 27 117
rect 33 111 39 117
rect 45 111 51 117
rect 57 111 63 117
rect 69 111 75 117
rect 81 111 87 117
rect 93 111 99 117
rect 105 111 111 117
rect 117 111 123 117
rect 129 111 135 117
rect 141 111 147 117
rect 153 111 159 117
rect 165 111 168 117
rect -36 108 168 111
<< mvnsubdiff >>
rect -36 357 168 360
rect -36 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 168 357
rect -36 348 168 351
rect -36 261 168 264
rect -36 255 -33 261
rect -27 255 -21 261
rect -15 255 -9 261
rect -3 255 3 261
rect 9 255 15 261
rect 21 255 27 261
rect 33 255 39 261
rect 45 255 51 261
rect 57 255 63 261
rect 69 255 75 261
rect 81 255 87 261
rect 93 255 99 261
rect 105 255 111 261
rect 117 255 123 261
rect 129 255 135 261
rect 141 255 147 261
rect 153 255 159 261
rect 165 255 168 261
rect -36 252 168 255
<< psubdiffcont >>
rect -45 399 -39 405
rect -33 399 -27 405
rect -21 399 -15 405
rect -9 399 -3 405
rect 3 399 9 405
rect 15 399 21 405
rect 27 399 33 405
rect 39 399 45 405
rect 51 399 57 405
rect 63 399 69 405
rect 75 399 81 405
rect 87 399 93 405
rect 99 399 105 405
rect 111 399 117 405
rect 123 399 129 405
rect 135 399 141 405
rect 147 399 153 405
rect 159 399 165 405
rect 171 399 177 405
rect -45 231 -39 237
rect -33 231 -27 237
rect -21 231 -15 237
rect -9 231 -3 237
rect 3 231 9 237
rect 15 231 21 237
rect 27 231 33 237
rect 39 231 45 237
rect 51 231 57 237
rect 63 231 69 237
rect 75 231 81 237
rect 87 231 93 237
rect 99 231 105 237
rect 111 231 117 237
rect 123 231 129 237
rect 135 231 141 237
rect 147 231 153 237
rect 159 231 165 237
rect 171 231 177 237
rect -45 39 -39 45
rect -33 39 -27 45
rect -21 39 -15 45
rect -9 39 -3 45
rect 3 39 9 45
rect 15 39 21 45
rect 27 39 33 45
rect 39 39 45 45
rect 51 39 57 45
rect 63 39 69 45
rect 75 39 81 45
rect 87 39 93 45
rect 99 39 105 45
rect 111 39 117 45
rect 123 39 129 45
rect 135 39 141 45
rect 147 39 153 45
rect 159 39 165 45
rect 171 39 177 45
rect -45 -33 -39 -27
rect -33 -33 -27 -27
rect -21 -33 -15 -27
rect -9 -33 -3 -27
rect 3 -33 9 -27
rect 15 -33 21 -27
rect 27 -33 33 -27
rect 39 -33 45 -27
rect 51 -33 57 -27
rect 63 -33 69 -27
rect 75 -33 81 -27
rect 87 -33 93 -27
rect 99 -33 105 -27
rect 111 -33 117 -27
rect 123 -33 129 -27
rect 135 -33 141 -27
rect 147 -33 153 -27
rect 159 -33 165 -27
rect 171 -33 177 -27
rect -45 -129 -39 -123
rect -33 -129 -27 -123
rect -21 -129 -15 -123
rect -9 -129 -3 -123
rect 3 -129 9 -123
rect 15 -129 21 -123
rect 27 -129 33 -123
rect 39 -129 45 -123
rect 51 -129 57 -123
rect 63 -129 69 -123
rect 75 -129 81 -123
rect 87 -129 93 -123
rect 99 -129 105 -123
rect 111 -129 117 -123
rect 123 -129 129 -123
rect 135 -129 141 -123
rect 147 -129 153 -123
rect 159 -129 165 -123
rect 171 -129 177 -123
<< nsubdiffcont >>
rect -33 207 -27 213
rect -21 207 -15 213
rect -9 207 -3 213
rect 3 207 9 213
rect 15 207 21 213
rect 27 207 33 213
rect 39 207 45 213
rect 51 207 57 213
rect 63 207 69 213
rect 75 207 81 213
rect 87 207 93 213
rect 99 207 105 213
rect 111 207 117 213
rect 123 207 129 213
rect 135 207 141 213
rect 147 207 153 213
rect 159 207 165 213
rect -33 111 -27 117
rect -21 111 -15 117
rect -9 111 -3 117
rect 3 111 9 117
rect 15 111 21 117
rect 27 111 33 117
rect 39 111 45 117
rect 51 111 57 117
rect 63 111 69 117
rect 75 111 81 117
rect 87 111 93 117
rect 99 111 105 117
rect 111 111 117 117
rect 123 111 129 117
rect 135 111 141 117
rect 147 111 153 117
rect 159 111 165 117
<< mvnsubdiffcont >>
rect -33 351 -27 357
rect -21 351 -15 357
rect -9 351 -3 357
rect 3 351 9 357
rect 15 351 21 357
rect 27 351 33 357
rect 39 351 45 357
rect 51 351 57 357
rect 63 351 69 357
rect 75 351 81 357
rect 87 351 93 357
rect 99 351 105 357
rect 111 351 117 357
rect 123 351 129 357
rect 135 351 141 357
rect 147 351 153 357
rect 159 351 165 357
rect -33 255 -27 261
rect -21 255 -15 261
rect -9 255 -3 261
rect 3 255 9 261
rect 15 255 21 261
rect 27 255 33 261
rect 39 255 45 261
rect 51 255 57 261
rect 63 255 69 261
rect 75 255 81 261
rect 87 255 93 261
rect 99 255 105 261
rect 111 255 117 261
rect 123 255 129 261
rect 135 255 141 261
rect 147 255 153 261
rect 159 255 165 261
<< polysilicon >>
rect -24 336 -12 342
rect 0 336 12 342
rect 24 336 36 342
rect 48 336 60 342
rect 72 336 84 342
rect 96 336 108 342
rect 120 336 132 342
rect 144 336 156 342
rect -24 288 -12 300
rect 0 288 12 300
rect 24 288 36 300
rect 48 288 60 300
rect -24 285 60 288
rect -24 279 -21 285
rect -15 279 -9 285
rect -3 279 3 285
rect 9 279 15 285
rect 21 279 27 285
rect 33 279 39 285
rect 45 279 51 285
rect 57 279 60 285
rect -24 276 60 279
rect 72 288 84 300
rect 96 288 108 300
rect 120 288 132 300
rect 144 288 156 300
rect 72 285 156 288
rect 72 279 75 285
rect 81 279 87 285
rect 93 279 99 285
rect 105 279 111 285
rect 117 279 123 285
rect 129 279 135 285
rect 141 279 147 285
rect 153 279 156 285
rect 72 276 156 279
rect -24 186 -12 192
rect 0 186 12 192
rect 24 186 36 192
rect 48 186 60 192
rect 72 186 84 192
rect 96 186 108 192
rect 120 186 132 192
rect 144 186 156 192
rect -24 144 -12 156
rect 0 144 12 156
rect 24 144 36 156
rect 48 144 60 156
rect 72 144 84 156
rect 96 144 108 156
rect 120 144 132 156
rect 144 144 156 156
rect -24 141 156 144
rect -24 135 -21 141
rect -15 135 -9 141
rect -3 135 3 141
rect 9 135 15 141
rect 21 135 27 141
rect 33 135 39 141
rect 45 135 51 141
rect 57 135 63 141
rect 69 135 75 141
rect 81 135 87 141
rect 93 135 99 141
rect 105 135 111 141
rect 117 135 123 141
rect 129 135 135 141
rect 141 135 147 141
rect 153 135 156 141
rect -24 132 156 135
rect -24 -51 156 -48
rect -24 -57 -21 -51
rect -15 -57 -9 -51
rect -3 -57 3 -51
rect 9 -57 15 -51
rect 21 -57 27 -51
rect 33 -57 39 -51
rect 45 -57 51 -51
rect 57 -57 63 -51
rect 69 -57 75 -51
rect 81 -57 87 -51
rect 93 -57 99 -51
rect 105 -57 111 -51
rect 117 -57 123 -51
rect 129 -57 135 -51
rect 141 -57 147 -51
rect 153 -57 156 -51
rect -24 -60 156 -57
rect -24 -72 -12 -60
rect 0 -72 12 -60
rect 24 -72 36 -60
rect 48 -72 60 -60
rect 72 -72 84 -60
rect 96 -72 108 -60
rect 120 -72 132 -60
rect 144 -72 156 -60
rect -24 -114 -12 -108
rect 0 -114 12 -108
rect 24 -114 36 -108
rect 48 -114 60 -108
rect 72 -114 84 -108
rect 96 -114 108 -108
rect 120 -114 132 -108
rect 144 -114 156 -108
<< polycontact >>
rect -21 279 -15 285
rect -9 279 -3 285
rect 3 279 9 285
rect 15 279 21 285
rect 27 279 33 285
rect 39 279 45 285
rect 51 279 57 285
rect 75 279 81 285
rect 87 279 93 285
rect 99 279 105 285
rect 111 279 117 285
rect 123 279 129 285
rect 135 279 141 285
rect 147 279 153 285
rect -21 135 -15 141
rect -9 135 -3 141
rect 3 135 9 141
rect 15 135 21 141
rect 27 135 33 141
rect 39 135 45 141
rect 51 135 57 141
rect 63 135 69 141
rect 75 135 81 141
rect 87 135 93 141
rect 99 135 105 141
rect 111 135 117 141
rect 123 135 129 141
rect 135 135 141 141
rect 147 135 153 141
rect -21 -57 -15 -51
rect -9 -57 -3 -51
rect 3 -57 9 -51
rect 15 -57 21 -51
rect 27 -57 33 -51
rect 39 -57 45 -51
rect 51 -57 57 -51
rect 63 -57 69 -51
rect 75 -57 81 -51
rect 87 -57 93 -51
rect 99 -57 105 -51
rect 111 -57 117 -51
rect 123 -57 129 -51
rect 135 -57 141 -51
rect 147 -57 153 -51
<< metal1 >>
rect -48 405 180 408
rect -48 399 -45 405
rect -39 399 -33 405
rect -27 399 -21 405
rect -15 399 -9 405
rect -3 399 3 405
rect 9 399 15 405
rect 21 399 27 405
rect 33 399 39 405
rect 45 399 51 405
rect 57 399 63 405
rect 69 399 75 405
rect 81 399 87 405
rect 93 399 99 405
rect 105 399 111 405
rect 117 399 123 405
rect 129 399 135 405
rect 141 399 147 405
rect 153 399 159 405
rect 165 399 171 405
rect 177 399 180 405
rect -48 396 180 399
rect -36 357 168 360
rect -36 351 -33 357
rect -27 351 -21 357
rect -15 351 -9 357
rect -3 351 3 357
rect 9 351 15 357
rect 21 351 27 357
rect 33 351 39 357
rect 45 351 51 357
rect 57 351 63 357
rect 69 351 75 357
rect 81 351 87 357
rect 93 351 99 357
rect 105 351 111 357
rect 117 351 123 357
rect 129 351 135 357
rect 141 351 147 357
rect 153 351 159 357
rect 165 351 168 357
rect -36 348 168 351
rect -36 333 -24 336
rect -36 327 -33 333
rect -27 327 -24 333
rect -36 321 -24 327
rect -36 315 -33 321
rect -27 315 -24 321
rect -36 309 -24 315
rect -36 303 -33 309
rect -27 303 -24 309
rect -36 300 -24 303
rect -12 333 0 336
rect -12 327 -9 333
rect -3 327 0 333
rect -12 321 0 327
rect -12 315 -9 321
rect -3 315 0 321
rect -12 309 0 315
rect -12 303 -9 309
rect -3 303 0 309
rect -12 300 0 303
rect 12 333 24 336
rect 12 327 15 333
rect 21 327 24 333
rect 12 321 24 327
rect 12 315 15 321
rect 21 315 24 321
rect 12 309 24 315
rect 12 303 15 309
rect 21 303 24 309
rect 12 300 24 303
rect 36 333 48 336
rect 36 327 39 333
rect 45 327 48 333
rect 36 321 48 327
rect 36 315 39 321
rect 45 315 48 321
rect 36 309 48 315
rect 36 303 39 309
rect 45 303 48 309
rect 36 300 48 303
rect 60 333 72 336
rect 60 327 63 333
rect 69 327 72 333
rect 60 321 72 327
rect 60 315 63 321
rect 69 315 72 321
rect 60 309 72 315
rect 60 303 63 309
rect 69 303 72 309
rect 60 300 72 303
rect 84 333 96 336
rect 84 327 87 333
rect 93 327 96 333
rect 84 321 96 327
rect 84 315 87 321
rect 93 315 96 321
rect 84 309 96 315
rect 84 303 87 309
rect 93 303 96 309
rect 84 300 96 303
rect 108 333 120 336
rect 108 327 111 333
rect 117 327 120 333
rect 108 321 120 327
rect 108 315 111 321
rect 117 315 120 321
rect 108 309 120 315
rect 108 303 111 309
rect 117 303 120 309
rect 108 300 120 303
rect 132 333 144 336
rect 132 327 135 333
rect 141 327 144 333
rect 132 321 144 327
rect 132 315 135 321
rect 141 315 144 321
rect 132 309 144 315
rect 132 303 135 309
rect 141 303 144 309
rect 132 300 144 303
rect 156 333 168 336
rect 156 327 159 333
rect 165 327 168 333
rect 156 321 168 327
rect 156 315 159 321
rect 165 315 168 321
rect 156 309 168 315
rect 156 303 159 309
rect 165 303 168 309
rect 156 300 168 303
rect -24 285 156 288
rect -24 279 -21 285
rect -15 279 -9 285
rect -3 279 3 285
rect 9 279 15 285
rect 21 279 27 285
rect 33 279 39 285
rect 45 279 51 285
rect 57 279 63 285
rect 69 279 75 285
rect 81 279 87 285
rect 93 279 99 285
rect 105 279 111 285
rect 117 279 123 285
rect 129 279 135 285
rect 141 279 147 285
rect 153 279 156 285
rect -24 276 156 279
rect -36 261 168 264
rect -36 255 -33 261
rect -27 255 -21 261
rect -15 255 -9 261
rect -3 255 3 261
rect 9 255 15 261
rect 21 255 27 261
rect 33 255 39 261
rect 45 255 51 261
rect 57 255 63 261
rect 69 255 75 261
rect 81 255 87 261
rect 93 255 99 261
rect 105 255 111 261
rect 117 255 123 261
rect 129 255 135 261
rect 141 255 147 261
rect 153 255 159 261
rect 165 255 168 261
rect -36 252 168 255
rect -48 237 180 240
rect -48 231 -45 237
rect -39 231 -33 237
rect -27 231 -21 237
rect -15 231 -9 237
rect -3 231 3 237
rect 9 231 15 237
rect 21 231 27 237
rect 33 231 39 237
rect 45 231 51 237
rect 57 231 63 237
rect 69 231 75 237
rect 81 231 87 237
rect 93 231 99 237
rect 105 231 111 237
rect 117 231 123 237
rect 129 231 135 237
rect 141 231 147 237
rect 153 231 159 237
rect 165 231 171 237
rect 177 231 180 237
rect -48 228 180 231
rect -48 213 180 216
rect -48 207 -33 213
rect -27 207 -21 213
rect -15 207 -9 213
rect -3 207 3 213
rect 9 207 15 213
rect 21 207 27 213
rect 33 207 39 213
rect 45 207 51 213
rect 57 207 63 213
rect 69 207 75 213
rect 81 207 87 213
rect 93 207 99 213
rect 105 207 111 213
rect 117 207 123 213
rect 129 207 135 213
rect 141 207 147 213
rect 153 207 159 213
rect 165 207 180 213
rect -48 204 180 207
rect -36 177 -24 186
rect -36 171 -33 177
rect -27 171 -24 177
rect -36 165 -24 171
rect -36 159 -33 165
rect -27 159 -24 165
rect -36 156 -24 159
rect -12 177 0 186
rect -12 171 -9 177
rect -3 171 0 177
rect -12 165 0 171
rect -12 159 -9 165
rect -3 159 0 165
rect -12 156 0 159
rect 12 177 24 186
rect 12 171 15 177
rect 21 171 24 177
rect 12 165 24 171
rect 12 159 15 165
rect 21 159 24 165
rect 12 156 24 159
rect 36 177 48 186
rect 36 171 39 177
rect 45 171 48 177
rect 36 165 48 171
rect 36 159 39 165
rect 45 159 48 165
rect 36 156 48 159
rect 60 177 72 186
rect 60 171 63 177
rect 69 171 72 177
rect 60 165 72 171
rect 60 159 63 165
rect 69 159 72 165
rect 60 156 72 159
rect 84 177 96 186
rect 84 171 87 177
rect 93 171 96 177
rect 84 165 96 171
rect 84 159 87 165
rect 93 159 96 165
rect 84 156 96 159
rect 108 177 120 186
rect 108 171 111 177
rect 117 171 120 177
rect 108 165 120 171
rect 108 159 111 165
rect 117 159 120 165
rect 108 156 120 159
rect 132 177 144 186
rect 132 171 135 177
rect 141 171 144 177
rect 132 165 144 171
rect 132 159 135 165
rect 141 159 144 165
rect 132 156 144 159
rect 156 177 168 186
rect 156 171 159 177
rect 165 171 168 177
rect 156 165 168 171
rect 156 159 159 165
rect 165 159 168 165
rect 156 156 168 159
rect -24 141 156 144
rect -24 135 -21 141
rect -15 135 -9 141
rect -3 135 3 141
rect 9 135 15 141
rect 21 135 27 141
rect 33 135 39 141
rect 45 135 51 141
rect 57 135 63 141
rect 69 135 75 141
rect 81 135 87 141
rect 93 135 99 141
rect 105 135 111 141
rect 117 135 123 141
rect 129 135 135 141
rect 141 135 147 141
rect 153 135 156 141
rect -24 132 156 135
rect -36 117 168 120
rect -36 111 -33 117
rect -27 111 -21 117
rect -15 111 -9 117
rect -3 111 3 117
rect 9 111 15 117
rect 21 111 27 117
rect 33 111 39 117
rect 45 111 51 117
rect 57 111 63 117
rect 69 111 75 117
rect 81 111 87 117
rect 93 111 99 117
rect 105 111 111 117
rect 117 111 123 117
rect 129 111 135 117
rect 141 111 147 117
rect 153 111 159 117
rect 165 111 168 117
rect -36 108 168 111
rect -48 45 180 48
rect -48 39 -45 45
rect -39 39 -33 45
rect -27 39 -21 45
rect -15 39 -9 45
rect -3 39 3 45
rect 9 39 15 45
rect 21 39 27 45
rect 33 39 39 45
rect 45 39 51 45
rect 57 39 63 45
rect 69 39 75 45
rect 81 39 87 45
rect 93 39 99 45
rect 105 39 111 45
rect 117 39 123 45
rect 129 39 135 45
rect 141 39 147 45
rect 153 39 159 45
rect 165 39 171 45
rect 177 39 180 45
rect -48 36 180 39
rect -48 -27 180 -24
rect -48 -33 -45 -27
rect -39 -33 -33 -27
rect -27 -33 -21 -27
rect -15 -33 -9 -27
rect -3 -33 3 -27
rect 9 -33 15 -27
rect 21 -33 27 -27
rect 33 -33 39 -27
rect 45 -33 51 -27
rect 57 -33 63 -27
rect 69 -33 75 -27
rect 81 -33 87 -27
rect 93 -33 99 -27
rect 105 -33 111 -27
rect 117 -33 123 -27
rect 129 -33 135 -27
rect 141 -33 147 -27
rect 153 -33 159 -27
rect 165 -33 171 -27
rect 177 -33 180 -27
rect -48 -36 180 -33
rect -24 -51 156 -48
rect -24 -57 -21 -51
rect -15 -57 -9 -51
rect -3 -57 3 -51
rect 9 -57 15 -51
rect 21 -57 27 -51
rect 33 -57 39 -51
rect 45 -57 51 -51
rect 57 -57 63 -51
rect 69 -57 75 -51
rect 81 -57 87 -51
rect 93 -57 99 -51
rect 105 -57 111 -51
rect 117 -57 123 -51
rect 129 -57 135 -51
rect 141 -57 147 -51
rect 153 -57 156 -51
rect -24 -60 156 -57
rect -36 -75 -24 -72
rect -36 -81 -33 -75
rect -27 -81 -24 -75
rect -36 -87 -24 -81
rect -36 -93 -33 -87
rect -27 -93 -24 -87
rect -36 -99 -24 -93
rect -36 -105 -33 -99
rect -27 -105 -24 -99
rect -36 -108 -24 -105
rect -12 -75 0 -72
rect -12 -81 -9 -75
rect -3 -81 0 -75
rect -12 -87 0 -81
rect -12 -93 -9 -87
rect -3 -93 0 -87
rect -12 -99 0 -93
rect -12 -105 -9 -99
rect -3 -105 0 -99
rect -12 -108 0 -105
rect 12 -75 24 -72
rect 12 -81 15 -75
rect 21 -81 24 -75
rect 12 -87 24 -81
rect 12 -93 15 -87
rect 21 -93 24 -87
rect 12 -99 24 -93
rect 12 -105 15 -99
rect 21 -105 24 -99
rect 12 -108 24 -105
rect 36 -75 48 -72
rect 36 -81 39 -75
rect 45 -81 48 -75
rect 36 -87 48 -81
rect 36 -93 39 -87
rect 45 -93 48 -87
rect 36 -99 48 -93
rect 36 -105 39 -99
rect 45 -105 48 -99
rect 36 -108 48 -105
rect 60 -75 72 -72
rect 60 -81 63 -75
rect 69 -81 72 -75
rect 60 -87 72 -81
rect 60 -93 63 -87
rect 69 -93 72 -87
rect 60 -99 72 -93
rect 60 -105 63 -99
rect 69 -105 72 -99
rect 60 -108 72 -105
rect 84 -75 96 -72
rect 84 -81 87 -75
rect 93 -81 96 -75
rect 84 -87 96 -81
rect 84 -93 87 -87
rect 93 -93 96 -87
rect 84 -99 96 -93
rect 84 -105 87 -99
rect 93 -105 96 -99
rect 84 -108 96 -105
rect 108 -75 120 -72
rect 108 -81 111 -75
rect 117 -81 120 -75
rect 108 -87 120 -81
rect 108 -93 111 -87
rect 117 -93 120 -87
rect 108 -99 120 -93
rect 108 -105 111 -99
rect 117 -105 120 -99
rect 108 -108 120 -105
rect 132 -75 144 -72
rect 132 -81 135 -75
rect 141 -81 144 -75
rect 132 -87 144 -81
rect 132 -93 135 -87
rect 141 -93 144 -87
rect 132 -99 144 -93
rect 132 -105 135 -99
rect 141 -105 144 -99
rect 132 -108 144 -105
rect 156 -75 168 -72
rect 156 -81 159 -75
rect 165 -81 168 -75
rect 156 -87 168 -81
rect 156 -93 159 -87
rect 165 -93 168 -87
rect 156 -99 168 -93
rect 156 -105 159 -99
rect 165 -105 168 -99
rect 156 -108 168 -105
rect -48 -123 180 -120
rect -48 -129 -45 -123
rect -39 -129 -33 -123
rect -27 -129 -21 -123
rect -15 -129 -9 -123
rect -3 -129 3 -123
rect 9 -129 15 -123
rect 21 -129 27 -123
rect 33 -129 39 -123
rect 45 -129 51 -123
rect 57 -129 63 -123
rect 69 -129 75 -123
rect 81 -129 87 -123
rect 93 -129 99 -123
rect 105 -129 111 -123
rect 117 -129 123 -123
rect 129 -129 135 -123
rect 141 -129 147 -123
rect 153 -129 159 -123
rect 165 -129 171 -123
rect 177 -129 180 -123
rect -48 -132 180 -129
<< via1 >>
rect -33 351 -27 357
rect 15 351 21 357
rect 63 351 69 357
rect 111 351 117 357
rect -33 327 -27 333
rect -33 315 -27 321
rect -33 303 -27 309
rect -9 327 -3 333
rect -9 315 -3 321
rect -9 303 -3 309
rect 15 327 21 333
rect 15 315 21 321
rect 15 303 21 309
rect 39 327 45 333
rect 39 315 45 321
rect 39 303 45 309
rect 63 327 69 333
rect 63 315 69 321
rect 63 303 69 309
rect 87 327 93 333
rect 87 315 93 321
rect 87 303 93 309
rect 111 327 117 333
rect 111 315 117 321
rect 111 303 117 309
rect 135 327 141 333
rect 135 315 141 321
rect 135 303 141 309
rect 159 327 165 333
rect 159 315 165 321
rect 159 303 165 309
rect 63 279 69 285
rect -33 171 -27 177
rect -33 159 -27 165
rect -9 171 -3 177
rect -9 159 -3 165
rect 15 171 21 177
rect 15 159 21 165
rect 39 171 45 177
rect 39 159 45 165
rect 63 171 69 177
rect 63 159 69 165
rect 87 171 93 177
rect 87 159 93 165
rect 111 171 117 177
rect 111 159 117 165
rect 135 171 141 177
rect 135 159 141 165
rect 159 171 165 177
rect 159 159 165 165
rect 63 135 69 141
rect -33 39 -27 45
rect 159 39 165 45
rect -33 -33 -27 -27
rect 159 -33 165 -27
rect 63 -57 69 -51
rect -33 -81 -27 -75
rect -33 -93 -27 -87
rect -33 -105 -27 -99
rect -9 -81 -3 -75
rect -9 -93 -3 -87
rect -9 -105 -3 -99
rect 15 -81 21 -75
rect 15 -93 21 -87
rect 15 -105 21 -99
rect 39 -81 45 -75
rect 39 -93 45 -87
rect 39 -105 45 -99
rect 63 -81 69 -75
rect 63 -93 69 -87
rect 63 -105 69 -99
rect 87 -81 93 -75
rect 87 -93 93 -87
rect 87 -105 93 -99
rect 111 -81 117 -75
rect 111 -93 117 -87
rect 111 -105 117 -99
rect 135 -81 141 -75
rect 135 -93 141 -87
rect 135 -105 141 -99
rect 159 -81 165 -75
rect 159 -93 165 -87
rect 159 -105 165 -99
rect -33 -129 -27 -123
rect 159 -129 165 -123
<< metal2 >>
rect -36 405 -24 408
rect -36 399 -33 405
rect -27 399 -24 405
rect -36 381 -24 399
rect -36 375 -33 381
rect -27 375 -24 381
rect -36 357 -24 375
rect -36 351 -33 357
rect -27 351 -24 357
rect -36 333 -24 351
rect 12 381 24 384
rect 12 375 15 381
rect 21 375 24 381
rect 12 357 24 375
rect 12 351 15 357
rect 21 351 24 357
rect -36 327 -33 333
rect -27 327 -24 333
rect -36 321 -24 327
rect -36 315 -33 321
rect -27 315 -24 321
rect -36 309 -24 315
rect -36 303 -33 309
rect -27 303 -24 309
rect -36 300 -24 303
rect -12 333 0 336
rect -12 327 -9 333
rect -3 327 0 333
rect -12 321 0 327
rect -12 315 -9 321
rect -3 315 0 321
rect -12 309 0 315
rect -12 303 -9 309
rect -3 303 0 309
rect -36 261 -24 264
rect -36 255 -33 261
rect -27 255 -24 261
rect -36 213 -24 255
rect -36 207 -33 213
rect -27 207 -24 213
rect -36 189 -24 207
rect -12 261 0 303
rect 12 333 24 351
rect 60 381 72 384
rect 60 375 63 381
rect 69 375 72 381
rect 60 357 72 375
rect 60 351 63 357
rect 69 351 72 357
rect 12 327 15 333
rect 21 327 24 333
rect 12 321 24 327
rect 12 315 15 321
rect 21 315 24 321
rect 12 309 24 315
rect 12 303 15 309
rect 21 303 24 309
rect 12 300 24 303
rect 36 333 48 336
rect 36 327 39 333
rect 45 327 48 333
rect 36 321 48 327
rect 36 315 39 321
rect 45 315 48 321
rect 36 309 48 315
rect 36 303 39 309
rect 45 303 48 309
rect -12 255 -9 261
rect -3 255 0 261
rect -12 213 0 255
rect -12 207 -9 213
rect -3 207 0 213
rect -12 204 0 207
rect 12 261 24 264
rect 12 255 15 261
rect 21 255 24 261
rect 12 213 24 255
rect 12 207 15 213
rect 21 207 24 213
rect -36 183 -33 189
rect -27 183 -24 189
rect 12 189 24 207
rect 36 261 48 303
rect 60 333 72 351
rect 108 381 120 384
rect 108 375 111 381
rect 117 375 120 381
rect 108 357 120 375
rect 108 351 111 357
rect 117 351 120 357
rect 60 327 63 333
rect 69 327 72 333
rect 60 321 72 327
rect 60 315 63 321
rect 69 315 72 321
rect 60 309 72 315
rect 60 303 63 309
rect 69 303 72 309
rect 60 300 72 303
rect 84 333 96 336
rect 84 327 87 333
rect 93 327 96 333
rect 84 321 96 327
rect 84 315 87 321
rect 93 315 96 321
rect 84 309 96 315
rect 84 303 87 309
rect 93 303 96 309
rect 60 285 72 288
rect 60 279 63 285
rect 69 279 72 285
rect 60 276 72 279
rect 36 255 39 261
rect 45 255 48 261
rect 36 213 48 255
rect 84 261 96 303
rect 108 333 120 351
rect 156 381 168 384
rect 156 375 159 381
rect 165 375 168 381
rect 156 357 168 375
rect 156 351 159 357
rect 165 351 168 357
rect 108 327 111 333
rect 117 327 120 333
rect 108 321 120 327
rect 108 315 111 321
rect 117 315 120 321
rect 108 309 120 315
rect 108 303 111 309
rect 117 303 120 309
rect 108 300 120 303
rect 132 333 144 336
rect 132 327 135 333
rect 141 327 144 333
rect 132 321 144 327
rect 132 315 135 321
rect 141 315 144 321
rect 132 309 144 315
rect 132 303 135 309
rect 141 303 144 309
rect 84 255 87 261
rect 93 255 96 261
rect 60 228 72 240
rect 36 207 39 213
rect 45 207 48 213
rect 36 204 48 207
rect 60 213 72 216
rect 60 207 63 213
rect 69 207 72 213
rect -36 177 -24 183
rect -36 171 -33 177
rect -27 171 -24 177
rect -36 165 -24 171
rect -36 159 -33 165
rect -27 159 -24 165
rect -36 156 -24 159
rect -12 177 0 186
rect -12 171 -9 177
rect -3 171 0 177
rect -12 165 0 171
rect -12 159 -9 165
rect -3 159 0 165
rect -36 117 -24 120
rect -36 111 -33 117
rect -27 111 -24 117
rect -36 45 -24 111
rect -36 39 -33 45
rect -27 39 -24 45
rect -36 -27 -24 39
rect -12 12 0 159
rect 12 183 15 189
rect 21 183 24 189
rect 60 189 72 207
rect 84 213 96 255
rect 84 207 87 213
rect 93 207 96 213
rect 84 204 96 207
rect 108 261 120 264
rect 108 255 111 261
rect 117 255 120 261
rect 108 213 120 255
rect 108 207 111 213
rect 117 207 120 213
rect 12 177 24 183
rect 12 171 15 177
rect 21 171 24 177
rect 12 165 24 171
rect 12 159 15 165
rect 21 159 24 165
rect 12 156 24 159
rect 36 177 48 186
rect 36 171 39 177
rect 45 171 48 177
rect 36 165 48 171
rect 36 159 39 165
rect 45 159 48 165
rect 36 12 48 159
rect 60 183 63 189
rect 69 183 72 189
rect 108 189 120 207
rect 132 261 144 303
rect 156 333 168 351
rect 156 327 159 333
rect 165 327 168 333
rect 156 321 168 327
rect 156 315 159 321
rect 165 315 168 321
rect 156 309 168 315
rect 156 303 159 309
rect 165 303 168 309
rect 156 300 168 303
rect 132 255 135 261
rect 141 255 144 261
rect 132 213 144 255
rect 132 207 135 213
rect 141 207 144 213
rect 132 204 144 207
rect 156 261 168 264
rect 156 255 159 261
rect 165 255 168 261
rect 156 213 168 255
rect 156 207 159 213
rect 165 207 168 213
rect 60 177 72 183
rect 60 171 63 177
rect 69 171 72 177
rect 60 165 72 171
rect 60 159 63 165
rect 69 159 72 165
rect 60 156 72 159
rect 84 177 96 186
rect 84 171 87 177
rect 93 171 96 177
rect 84 165 96 171
rect 84 159 87 165
rect 93 159 96 165
rect 60 141 72 144
rect 60 135 63 141
rect 69 135 72 141
rect 60 132 72 135
rect -12 9 48 12
rect -12 3 -9 9
rect -3 3 15 9
rect 21 3 39 9
rect 45 3 48 9
rect -12 0 48 3
rect 84 12 96 159
rect 108 183 111 189
rect 117 183 120 189
rect 156 189 168 207
rect 108 177 120 183
rect 108 171 111 177
rect 117 171 120 177
rect 108 165 120 171
rect 108 159 111 165
rect 117 159 120 165
rect 108 156 120 159
rect 132 177 144 186
rect 132 171 135 177
rect 141 171 144 177
rect 132 165 144 171
rect 132 159 135 165
rect 141 159 144 165
rect 132 12 144 159
rect 156 183 159 189
rect 165 183 168 189
rect 156 177 168 183
rect 156 171 159 177
rect 165 171 168 177
rect 156 165 168 171
rect 156 159 159 165
rect 165 159 168 165
rect 156 156 168 159
rect 84 9 144 12
rect 84 3 87 9
rect 93 3 111 9
rect 117 3 135 9
rect 141 3 144 9
rect 84 0 144 3
rect 156 117 168 120
rect 156 111 159 117
rect 165 111 168 117
rect 156 45 168 111
rect 156 39 159 45
rect 165 39 168 45
rect -36 -33 -33 -27
rect -27 -33 -24 -27
rect -36 -75 -24 -33
rect -36 -81 -33 -75
rect -27 -81 -24 -75
rect -36 -87 -24 -81
rect -36 -93 -33 -87
rect -27 -93 -24 -87
rect -36 -99 -24 -93
rect -36 -105 -33 -99
rect -27 -105 -24 -99
rect -36 -123 -24 -105
rect -12 -75 0 -72
rect -12 -81 -9 -75
rect -3 -81 0 -75
rect -12 -87 0 -81
rect -12 -93 -9 -87
rect -3 -93 0 -87
rect -12 -99 0 -93
rect -12 -105 -9 -99
rect -3 -105 0 -99
rect -12 -108 0 -105
rect 12 -75 24 0
rect 60 -51 72 -48
rect 60 -57 63 -51
rect 69 -57 72 -51
rect 60 -60 72 -57
rect 12 -81 15 -75
rect 21 -81 24 -75
rect 12 -87 24 -81
rect 12 -93 15 -87
rect 21 -93 24 -87
rect 12 -99 24 -93
rect 12 -105 15 -99
rect 21 -105 24 -99
rect 12 -108 24 -105
rect 36 -75 48 -72
rect 36 -81 39 -75
rect 45 -81 48 -75
rect 36 -87 48 -81
rect 36 -93 39 -87
rect 45 -93 48 -87
rect 36 -99 48 -93
rect 36 -105 39 -99
rect 45 -105 48 -99
rect 36 -108 48 -105
rect 60 -75 72 -72
rect 60 -81 63 -75
rect 69 -81 72 -75
rect 60 -87 72 -81
rect 60 -93 63 -87
rect 69 -93 72 -87
rect 60 -99 72 -93
rect 60 -105 63 -99
rect 69 -105 72 -99
rect 60 -108 72 -105
rect 84 -75 96 -72
rect 84 -81 87 -75
rect 93 -81 96 -75
rect 84 -87 96 -81
rect 84 -93 87 -87
rect 93 -93 96 -87
rect 84 -99 96 -93
rect 84 -105 87 -99
rect 93 -105 96 -99
rect 84 -108 96 -105
rect 108 -75 120 0
rect 156 -27 168 39
rect 156 -33 159 -27
rect 165 -33 168 -27
rect 108 -81 111 -75
rect 117 -81 120 -75
rect 108 -87 120 -81
rect 108 -93 111 -87
rect 117 -93 120 -87
rect 108 -99 120 -93
rect 108 -105 111 -99
rect 117 -105 120 -99
rect 108 -108 120 -105
rect 132 -75 144 -72
rect 132 -81 135 -75
rect 141 -81 144 -75
rect 132 -87 144 -81
rect 132 -93 135 -87
rect 141 -93 144 -87
rect 132 -99 144 -93
rect 132 -105 135 -99
rect 141 -105 144 -99
rect 132 -108 144 -105
rect 156 -75 168 -33
rect 156 -81 159 -75
rect 165 -81 168 -75
rect 156 -87 168 -81
rect 156 -93 159 -87
rect 165 -93 168 -87
rect 156 -99 168 -93
rect 156 -105 159 -99
rect 165 -105 168 -99
rect -36 -129 -33 -123
rect -27 -129 -24 -123
rect -36 -132 -24 -129
rect 156 -123 168 -105
rect 156 -129 159 -123
rect 165 -129 168 -123
rect 156 -132 168 -129
<< via2 >>
rect -33 399 -27 405
rect -33 375 -27 381
rect -33 351 -27 357
rect 15 375 21 381
rect 15 351 21 357
rect -33 327 -27 333
rect -33 303 -27 309
rect -33 255 -27 261
rect -33 207 -27 213
rect 63 375 69 381
rect 63 351 69 357
rect 15 327 21 333
rect 15 303 21 309
rect -9 255 -3 261
rect -9 207 -3 213
rect 15 255 21 261
rect 15 207 21 213
rect -33 183 -27 189
rect 111 375 117 381
rect 111 351 117 357
rect 63 327 69 333
rect 63 303 69 309
rect 63 279 69 285
rect 39 255 45 261
rect 159 375 165 381
rect 159 351 165 357
rect 111 327 117 333
rect 111 303 117 309
rect 87 255 93 261
rect 39 207 45 213
rect 63 207 69 213
rect -33 159 -27 165
rect -33 111 -27 117
rect -33 39 -27 45
rect 15 183 21 189
rect 87 207 93 213
rect 111 255 117 261
rect 111 207 117 213
rect 15 159 21 165
rect 63 183 69 189
rect 159 327 165 333
rect 159 303 165 309
rect 135 255 141 261
rect 135 207 141 213
rect 159 255 165 261
rect 159 207 165 213
rect 63 159 69 165
rect 63 135 69 141
rect -9 3 -3 9
rect 15 3 21 9
rect 39 3 45 9
rect 111 183 117 189
rect 111 159 117 165
rect 159 183 165 189
rect 159 159 165 165
rect 87 3 93 9
rect 111 3 117 9
rect 135 3 141 9
rect 159 111 165 117
rect 159 39 165 45
rect -33 -33 -27 -27
rect -33 -81 -27 -75
rect -33 -105 -27 -99
rect 63 -57 69 -51
rect 63 -81 69 -75
rect 63 -105 69 -99
rect 159 -33 165 -27
rect 159 -81 165 -75
rect 159 -105 165 -99
rect -33 -129 -27 -123
rect 159 -129 165 -123
<< metal3 >>
rect -48 405 180 408
rect -48 399 -33 405
rect -27 399 180 405
rect -48 396 180 399
rect -48 381 180 384
rect -48 375 -33 381
rect -27 375 15 381
rect 21 375 63 381
rect 69 375 111 381
rect 117 375 159 381
rect 165 375 180 381
rect -48 372 180 375
rect -48 357 180 360
rect -48 351 -33 357
rect -27 351 15 357
rect 21 351 63 357
rect 69 351 111 357
rect 117 351 159 357
rect 165 351 180 357
rect -48 333 180 351
rect -48 327 -33 333
rect -27 327 15 333
rect 21 327 63 333
rect 69 327 111 333
rect 117 327 159 333
rect 165 327 180 333
rect -48 309 180 327
rect -48 303 -33 309
rect -27 303 15 309
rect 21 303 63 309
rect 69 303 111 309
rect 117 303 159 309
rect 165 303 180 309
rect -48 300 180 303
rect 60 285 72 288
rect 60 279 63 285
rect 69 279 72 285
rect 60 276 72 279
rect -48 261 180 264
rect -48 255 -33 261
rect -27 255 -9 261
rect -3 255 15 261
rect 21 255 39 261
rect 45 255 87 261
rect 93 255 111 261
rect 117 255 135 261
rect 141 255 159 261
rect 165 255 180 261
rect -48 246 180 255
rect -48 237 180 240
rect -48 231 63 237
rect 69 231 180 237
rect -48 228 180 231
rect -48 213 180 222
rect -48 207 -33 213
rect -27 207 -9 213
rect -3 207 15 213
rect 21 207 39 213
rect 45 207 63 213
rect 69 207 87 213
rect 93 207 111 213
rect 117 207 135 213
rect 141 207 159 213
rect 165 207 180 213
rect -48 204 180 207
rect -48 189 180 192
rect -48 183 -33 189
rect -27 183 15 189
rect 21 183 63 189
rect 69 183 111 189
rect 117 183 159 189
rect 165 183 180 189
rect -48 180 180 183
rect -48 165 180 168
rect -48 159 -33 165
rect -27 159 15 165
rect 21 159 63 165
rect 69 159 111 165
rect 117 159 159 165
rect 165 159 180 165
rect -48 156 180 159
rect 60 141 72 144
rect 60 135 63 141
rect 69 135 72 141
rect 60 132 72 135
rect -48 117 168 120
rect -48 111 -33 117
rect -27 111 159 117
rect 165 111 168 117
rect -48 108 168 111
rect -48 81 180 96
rect -48 75 63 81
rect 69 75 180 81
rect -48 60 180 75
rect -48 45 180 48
rect -48 39 -33 45
rect -27 39 159 45
rect 165 39 180 45
rect -48 36 180 39
rect -48 9 180 24
rect -48 3 -9 9
rect -3 3 15 9
rect 21 3 39 9
rect 45 3 87 9
rect 93 3 111 9
rect 117 3 135 9
rect 141 3 180 9
rect -48 -12 180 3
rect -48 -27 180 -24
rect -48 -33 -33 -27
rect -27 -33 159 -27
rect 165 -33 180 -27
rect -48 -36 180 -33
rect 60 -51 72 -48
rect 60 -57 63 -51
rect 69 -57 72 -51
rect 60 -60 72 -57
rect -48 -75 180 -72
rect -48 -81 -33 -75
rect -27 -81 63 -75
rect 69 -81 159 -75
rect 165 -81 180 -75
rect -48 -99 180 -81
rect -48 -105 -33 -99
rect -27 -105 63 -99
rect 69 -105 159 -99
rect 165 -105 180 -99
rect -48 -123 180 -105
rect -48 -129 -33 -123
rect -27 -129 159 -123
rect 165 -129 180 -123
rect -48 -132 180 -129
<< via3 >>
rect 63 279 69 285
rect -33 255 -27 261
rect -9 255 -3 261
rect 15 255 21 261
rect 39 255 45 261
rect 87 255 93 261
rect 111 255 117 261
rect 135 255 141 261
rect 159 255 165 261
rect 63 231 69 237
rect -33 207 -27 213
rect -9 207 -3 213
rect 15 207 21 213
rect 39 207 45 213
rect 63 207 69 213
rect 87 207 93 213
rect 111 207 117 213
rect 135 207 141 213
rect 159 207 165 213
rect 63 135 69 141
rect 63 75 69 81
rect 63 -57 69 -51
<< metal4 >>
rect 60 285 72 288
rect 60 279 63 285
rect 69 279 72 285
rect -36 261 -24 264
rect -36 255 -33 261
rect -27 255 -24 261
rect -36 213 -24 255
rect -36 207 -33 213
rect -27 207 -24 213
rect -36 204 -24 207
rect -12 261 0 264
rect -12 255 -9 261
rect -3 255 0 261
rect -12 213 0 255
rect -12 207 -9 213
rect -3 207 0 213
rect -12 204 0 207
rect 12 261 24 264
rect 12 255 15 261
rect 21 255 24 261
rect 12 213 24 255
rect 12 207 15 213
rect 21 207 24 213
rect 12 204 24 207
rect 36 261 48 264
rect 36 255 39 261
rect 45 255 48 261
rect 36 213 48 255
rect 60 237 72 279
rect 60 231 63 237
rect 69 231 72 237
rect 60 228 72 231
rect 84 261 96 264
rect 84 255 87 261
rect 93 255 96 261
rect 36 207 39 213
rect 45 207 48 213
rect 36 204 48 207
rect 60 213 72 216
rect 60 207 63 213
rect 69 207 72 213
rect 60 204 72 207
rect 84 213 96 255
rect 84 207 87 213
rect 93 207 96 213
rect 84 204 96 207
rect 108 261 120 264
rect 108 255 111 261
rect 117 255 120 261
rect 108 213 120 255
rect 108 207 111 213
rect 117 207 120 213
rect 108 204 120 207
rect 132 261 144 264
rect 132 255 135 261
rect 141 255 144 261
rect 132 213 144 255
rect 132 207 135 213
rect 141 207 144 213
rect 132 204 144 207
rect 156 261 168 264
rect 156 255 159 261
rect 165 255 168 261
rect 156 213 168 255
rect 156 207 159 213
rect 165 207 168 213
rect 156 204 168 207
rect 60 141 72 144
rect 60 135 63 141
rect 69 135 72 141
rect 60 81 72 135
rect 60 75 63 81
rect 69 75 72 81
rect 60 -51 72 75
rect 60 -57 63 -51
rect 69 -57 72 -51
rect 60 -60 72 -57
<< labels >>
rlabel metal3 -48 -132 180 -120 0 vss
port 7 nsew
rlabel metal3 -48 0 180 12 0 out
port 2 nsew
rlabel metal3 -48 72 180 84 0 in
port 1 nsew
rlabel metal3 -48 228 180 240 0 gp
port 4 nsew
rlabel metal1 -48 204 180 216 0 bp
port 6 nsew
rlabel metal3 -48 252 -36 264 0 vdx
port 5 nsew
rlabel metal3 -48 372 180 384 0 vdh
port 3 nsew
rlabel metal2 -12 -96 0 -84 0 d1
rlabel metal2 36 -96 48 -84 0 d2
rlabel metal2 132 -96 144 -84 0 d4
rlabel metal2 84 -96 96 -84 0 d3
<< end >>
