magic
tech gf180mcuC
timestamp 1665149341
<< via2 >>
rect -780 228 -768 288
rect -60 228 -48 288
rect 60 228 72 288
rect 780 228 792 288
rect -540 132 -528 144
rect -420 132 -408 144
rect 420 132 432 144
rect 540 132 552 144
rect -300 84 -288 96
rect 300 84 312 96
rect -660 -60 -648 0
rect -180 -60 -168 0
rect 180 -60 192 0
rect 660 -60 672 0
<< metal3 >>
rect -936 528 -924 588
rect -936 480 -924 492
rect -936 456 -924 468
rect -936 324 -924 336
rect -936 228 -924 288
rect -936 180 -924 192
rect -936 132 -924 144
rect -936 84 -924 96
rect -936 36 -924 48
rect -936 -60 -924 0
rect -936 -180 -924 -120
<< via3 >>
rect -396 228 -384 288
rect 396 228 408 288
rect -804 180 -792 192
rect -36 180 -24 192
rect 36 180 48 192
rect 804 180 816 192
rect -516 132 -504 144
rect -444 132 -432 144
rect -324 132 -312 144
rect 324 132 336 144
rect 444 132 456 144
rect 516 132 528 144
rect -756 84 -744 96
rect -684 84 -672 96
rect -276 84 -264 96
rect -156 84 -144 96
rect -84 84 -72 96
rect 84 84 96 96
rect 156 84 168 96
rect 276 84 288 96
rect 684 84 696 96
rect 756 84 768 96
rect -636 36 -624 48
rect -204 36 -192 48
rect 204 36 216 48
rect 636 36 648 48
rect -564 -60 -552 0
rect 564 -60 576 0
use manf_cell  manf_cell_0
timestamp 1663176840
transform 1 0 -120 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_1
timestamp 1663176840
transform 1 0 0 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_2
timestamp 1663176840
transform 1 0 120 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_3
timestamp 1663176840
transform 1 0 240 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_4
timestamp 1663176840
transform 1 0 360 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_5
timestamp 1663176840
transform 1 0 480 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_6
timestamp 1663176840
transform 1 0 600 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_9
timestamp 1663176840
transform -1 0 132 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_10
timestamp 1663176840
transform -1 0 12 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_11
timestamp 1663176840
transform -1 0 -108 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_12
timestamp 1663176840
transform -1 0 -228 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_13
timestamp 1663176840
transform -1 0 -348 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_14
timestamp 1663176840
transform -1 0 -468 0 1 -48
box -720 -132 -588 660
use manf_cell  manf_cell_16
timestamp 1663176840
transform -1 0 -588 0 1 -48
box -720 -132 -588 660
use manf_edge  manf_edge_0
timestamp 1663179863
transform 1 0 -168 0 1 -48
box -756 -132 -660 660
use manf_edge  manf_edge_1
timestamp 1663179863
transform -1 0 180 0 1 -48
box -756 -132 -660 660
<< labels >>
rlabel metal3 -936 36 -924 48 0 ip
port 1 nsew
rlabel metal3 -936 180 -924 192 0 im
port 2 nsew
rlabel metal3 -936 228 -924 288 0 op
port 3 nsew
rlabel metal3 -936 -60 -924 0 0 om
port 4 nsew
rlabel metal3 -936 528 -924 588 0 vdd
port 5 nsew
rlabel metal3 -936 456 -924 468 0 gp
port 6 nsew
rlabel metal3 -936 324 -924 336 0 bp
port 7 nsew
rlabel metal3 -936 480 -924 492 0 vreg
port 8 nsew
rlabel metal3 -936 -180 -924 -120 0 gnd
port 9 nsew
rlabel metal3 -936 132 -924 144 0 x
rlabel metal3 -936 84 -924 96 0 y
<< end >>
