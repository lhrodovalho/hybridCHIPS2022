magic
tech gf180mcuC
timestamp 1665134701
<< via2 >>
rect -768 324 -756 348
rect -648 324 -636 348
rect 792 324 804 348
rect 912 324 924 348
rect 1272 324 1284 348
rect 1392 324 1404 348
rect 2832 324 2844 348
rect 2952 324 2964 348
rect -288 300 -276 312
rect 432 300 444 312
rect 1752 300 1764 312
rect 2472 300 2484 312
rect -768 264 -756 288
rect -648 264 -636 288
rect 792 264 804 288
rect 912 264 924 288
rect 1272 264 1284 288
rect 1392 264 1404 288
rect 2832 264 2844 288
rect 2952 264 2964 288
rect -168 168 -156 180
rect 312 168 324 180
rect 1872 168 1884 180
rect 2352 168 2364 180
rect -48 120 -36 132
rect 72 120 84 132
rect 192 120 204 132
rect 1992 120 2004 132
rect 2112 120 2124 132
rect 2232 120 2244 132
rect -888 12 -876 36
rect -528 12 -516 36
rect 672 12 684 36
rect 1032 12 1044 36
rect 1152 12 1164 36
rect 1512 12 1524 36
rect 2712 12 2724 36
rect 3072 12 3084 36
rect -408 -12 -396 0
rect 552 -12 564 0
rect 1632 -12 1644 0
rect 2592 -12 2604 0
rect -888 -48 -876 -24
rect -528 -48 -516 -24
rect 672 -48 684 -24
rect 1032 -48 1044 -24
rect 1152 -48 1164 -24
rect 1512 -48 1524 -24
rect 2712 -48 2724 -24
rect 3072 -48 3084 -24
<< mimcap >>
rect -1020 840 2976 888
rect -1020 756 -1008 840
rect -924 756 2976 840
rect -1020 744 2976 756
rect -1020 -252 2976 -240
rect -1020 -336 -1008 -252
rect -924 -336 2976 -252
rect -1020 -384 2976 -336
<< mimcapcontact >>
rect -1008 756 -924 840
rect -1008 -336 -924 -252
<< metal3 >>
rect -1044 588 -1032 648
rect -1044 534 -1032 552
rect -1044 516 -1032 528
rect -1044 384 -1032 396
rect -1104 346 -1032 348
rect -1104 320 -1102 346
rect -1094 320 -1054 346
rect -1046 320 -1032 346
rect -1104 318 -1032 320
rect -1104 310 -1032 312
rect -1104 302 -1078 310
rect -1070 302 -1032 310
rect -1104 300 -1032 302
rect -1104 292 -1032 294
rect -1104 266 -1102 292
rect -1094 266 -1054 292
rect -1046 266 -1032 292
rect -1104 264 -1032 266
rect -1044 216 -1032 228
rect -1044 168 -1032 180
rect -1044 120 -1032 132
rect -1044 72 -1032 84
rect -1104 34 -1032 36
rect -1104 8 -1102 34
rect -1094 8 -1054 34
rect -1046 8 -1032 34
rect -1104 6 -1032 8
rect -1104 -2 -1032 0
rect -1104 -10 -1078 -2
rect -1070 -10 -1032 -2
rect -1104 -12 -1032 -10
rect -1104 -20 -1032 -18
rect -1104 -46 -1102 -20
rect -1094 -46 -1054 -20
rect -1046 -46 -1032 -20
rect -1104 -48 -1032 -46
rect -1044 -168 -1032 -108
<< via3 >>
rect -1102 320 -1094 346
rect -1054 320 -1046 346
rect 168 324 180 348
rect 2016 324 2028 348
rect -1078 302 -1070 310
rect -744 300 -732 312
rect -672 300 -660 312
rect 336 300 348 312
rect 816 300 828 312
rect 888 300 900 312
rect 1296 300 1308 312
rect 1368 300 1380 312
rect 1848 300 1860 312
rect 2856 300 2868 312
rect 2928 300 2940 312
rect -1102 266 -1094 292
rect -1054 266 -1046 292
rect 168 264 180 288
rect 2016 264 2028 288
rect -792 216 -780 228
rect -624 216 -612 228
rect -432 216 -420 228
rect 576 216 588 228
rect 768 216 780 228
rect 936 216 948 228
rect 1248 216 1260 228
rect 1416 216 1428 228
rect 1608 216 1620 228
rect 2616 216 2628 228
rect 2808 216 2820 228
rect 2976 216 2988 228
rect -144 168 -132 180
rect -72 168 -60 180
rect 216 168 228 180
rect 288 168 300 180
rect 1896 168 1908 180
rect 1968 168 1980 180
rect 2256 168 2268 180
rect 2328 168 2340 180
rect -384 120 -372 132
rect -312 120 -300 132
rect 48 120 60 132
rect 96 120 108 132
rect 456 120 468 132
rect 528 120 540 132
rect 1656 120 1668 132
rect 1728 120 1740 132
rect 2088 120 2100 132
rect 2136 120 2148 132
rect 2496 120 2508 132
rect 2568 120 2580 132
rect -864 72 -852 84
rect -552 72 -540 84
rect -264 72 -252 84
rect 408 72 420 84
rect 696 72 708 84
rect 1008 72 1020 84
rect 1176 72 1188 84
rect 1488 72 1500 84
rect 1776 72 1788 84
rect 2448 72 2460 84
rect 2736 72 2748 84
rect 3048 72 3060 84
rect -1102 8 -1094 34
rect -1054 8 -1046 34
rect -24 12 -12 36
rect 2208 12 2220 36
rect -1078 -10 -1070 -2
rect -912 -12 -900 0
rect -504 -12 -492 0
rect -192 -12 -180 0
rect 648 -12 660 0
rect 1056 -12 1068 0
rect 1128 -12 1140 0
rect 1536 -12 1548 0
rect 2376 -12 2388 0
rect 2688 -12 2700 0
rect 3096 -12 3108 0
rect -1102 -46 -1094 -20
rect -1054 -46 -1046 -20
rect -24 -48 -12 -24
rect 2208 -48 2220 -24
<< metal4 >>
rect -1032 888 2988 900
rect -1104 744 -1092 756
rect -1104 696 -1092 732
rect -1104 346 -1092 684
rect -1104 320 -1102 346
rect -1094 320 -1092 346
rect -1104 292 -1092 320
rect -1104 266 -1102 292
rect -1094 266 -1092 292
rect -1104 264 -1092 266
rect -1080 720 -1068 756
rect -1080 310 -1068 708
rect -1080 302 -1078 310
rect -1070 302 -1068 310
rect -1080 264 -1068 302
rect -1056 744 -1044 756
rect -1056 696 -1044 732
rect -1032 744 -1020 888
rect 2976 744 2988 888
rect -1032 720 2988 744
rect -1032 708 -1020 720
rect 2976 708 2988 720
rect -1056 346 -1044 684
rect -1056 320 -1054 346
rect -1046 320 -1044 346
rect -1056 292 -1044 320
rect -1056 266 -1054 292
rect -1046 266 -1044 292
rect -1056 264 -1044 266
rect -1104 34 -1092 36
rect -1104 8 -1102 34
rect -1094 8 -1092 34
rect -1104 -20 -1092 8
rect -1104 -46 -1102 -20
rect -1094 -46 -1092 -20
rect -1104 -180 -1092 -46
rect -1104 -228 -1092 -192
rect -1104 -252 -1092 -240
rect -1080 -2 -1068 36
rect -1080 -10 -1078 -2
rect -1070 -10 -1068 -2
rect -1080 -204 -1068 -10
rect -1080 -252 -1068 -216
rect -1056 34 -1044 36
rect -1056 8 -1054 34
rect -1046 8 -1044 34
rect -1056 -20 -1044 8
rect -1056 -46 -1054 -20
rect -1046 -46 -1044 -20
rect -1056 -180 -1044 -46
rect -1056 -228 -1044 -192
rect -1056 -252 -1044 -240
rect -1032 -216 -1020 -204
rect 2976 -216 2988 -204
rect -1032 -240 2988 -216
rect -1032 -384 -1020 -240
rect 2976 -384 2988 -240
rect -1032 -396 2988 -384
<< via4 >>
rect -1104 732 -1092 744
rect -1104 684 -1092 696
rect -1080 708 -1068 720
rect -1056 732 -1044 744
rect -1020 708 2976 720
rect -1056 684 -1044 696
rect -1104 -192 -1092 -180
rect -1104 -240 -1092 -228
rect -1080 -216 -1068 -204
rect -1056 -192 -1044 -180
rect -1056 -240 -1044 -228
rect -1020 -216 2976 -204
<< metal5 >>
rect -1032 840 2988 900
rect -1032 756 -1008 840
rect -924 756 2988 840
rect -1032 744 2988 756
rect -1116 732 -1104 744
rect -1092 732 -1056 744
rect -1044 732 2988 744
rect -1116 708 -1080 720
rect -1068 708 -1020 720
rect 2976 708 2988 720
rect -1116 684 -1104 696
rect -1092 684 -1056 696
rect -1044 684 2988 696
rect -1116 -192 -1104 -180
rect -1092 -192 -1056 -180
rect -1044 -192 2988 -180
rect -1116 -216 -1080 -204
rect -1068 -216 -1020 -204
rect 2976 -216 2988 -204
rect -1116 -240 -1104 -228
rect -1092 -240 -1056 -228
rect -1044 -240 2988 -228
rect -1032 -252 2988 -240
rect -1032 -336 -1008 -252
rect -924 -336 2988 -252
rect -1032 -396 2988 -336
use manfvieru_cell  manfvieru_cell_0
timestamp 1664997892
transform 1 0 252 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_1
timestamp 1664997892
transform 1 0 372 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_2
timestamp 1664997892
transform 1 0 492 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_3
timestamp 1664997892
transform 1 0 612 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_4
timestamp 1664997892
transform 1 0 732 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_5
timestamp 1664997892
transform 1 0 852 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_6
timestamp 1664997892
transform 1 0 972 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_7
timestamp 1664997892
transform 1 0 1092 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_8
timestamp 1664997892
transform 1 0 1212 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_9
timestamp 1664997892
transform 1 0 1332 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_10
timestamp 1664997892
transform 1 0 1452 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_11
timestamp 1664997892
transform -1 0 264 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_12
timestamp 1664997892
transform -1 0 384 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_13
timestamp 1664997892
transform -1 0 -1176 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_14
timestamp 1664997892
transform 1 0 -228 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_15
timestamp 1664997892
transform -1 0 -1296 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_16
timestamp 1664997892
transform 1 0 -108 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_17
timestamp 1664997892
transform -1 0 2424 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_18
timestamp 1664997892
transform 1 0 3492 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_19
timestamp 1664997892
transform -1 0 2304 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_20
timestamp 1664997892
transform -1 0 1944 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_21
timestamp 1664997892
transform 1 0 3372 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_22
timestamp 1664997892
transform -1 0 1704 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_23
timestamp 1664997892
transform -1 0 1824 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_24
timestamp 1664997892
transform -1 0 1464 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_25
timestamp 1664997892
transform -1 0 1584 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_26
timestamp 1664997892
transform -1 0 1224 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_27
timestamp 1664997892
transform -1 0 1344 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_28
timestamp 1664997892
transform -1 0 1104 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_29
timestamp 1664997892
transform -1 0 984 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_30
timestamp 1664997892
transform -1 0 744 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_31
timestamp 1664997892
transform -1 0 864 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_32
timestamp 1664997892
transform 1 0 1812 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_33
timestamp 1664997892
transform 1 0 1932 0 1 -36
box -720 -132 -588 708
use manfvieru_edge  manfvieru_edge_0
timestamp 1664998004
transform 1 0 -276 0 1 -36
box -756 -132 -660 708
use manfvieru_edge  manfvieru_edge_1
timestamp 1664998004
transform -1 0 2472 0 1 -36
box -756 -132 -660 708
<< labels >>
rlabel metal3 -1044 -168 -1032 -108 0 gnd
port 9 nsew
rlabel metal3 -1044 -48 -1032 -36 0 om
port 4 nsew
rlabel metal3 -1044 -12 -1032 0 0 xp
rlabel metal3 -1044 588 -1032 648 0 vdd
port 5 nsew
rlabel metal3 -1044 516 -1032 528 0 gp
port 6 nsew
rlabel metal3 -1044 384 -1032 396 0 bp
port 7 nsew
rlabel metal3 -1044 540 -1032 552 0 vreg
port 8 nsew
rlabel metal3 -1044 216 -1032 228 0 im
port 2 nsew
rlabel metal3 -1044 336 -1032 348 0 op
port 3 nsew
rlabel metal3 -1044 300 -1032 312 0 xm
rlabel metal3 -1044 168 -1032 180 0 x
rlabel metal3 -1044 72 -1032 84 0 ip
port 1 nsew
rlabel metal3 -1044 120 -1032 132 0 y
<< end >>
