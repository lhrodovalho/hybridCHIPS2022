magic
tech gf180mcuC
timestamp 1664997892
<< nwell >>
rect -720 570 -588 690
rect -720 414 -588 546
<< nmos >>
rect -696 -108 -684 -72
rect -672 -108 -660 -72
rect -648 -108 -636 -72
rect -624 -108 -612 -72
<< pmos >>
rect -696 468 -684 498
rect -672 468 -660 498
rect -648 468 -636 498
rect -624 468 -612 498
<< mvpmos >>
rect -696 624 -684 660
rect -672 624 -660 660
rect -648 624 -636 660
rect -624 624 -612 660
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
<< pdiff >>
rect -708 489 -696 498
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 477 -696 483
rect -708 471 -705 477
rect -699 471 -696 477
rect -708 468 -696 471
rect -684 489 -672 498
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 477 -672 483
rect -684 471 -681 477
rect -675 471 -672 477
rect -684 468 -672 471
rect -660 489 -648 498
rect -660 483 -657 489
rect -651 483 -648 489
rect -660 477 -648 483
rect -660 471 -657 477
rect -651 471 -648 477
rect -660 468 -648 471
rect -636 489 -624 498
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 477 -624 483
rect -636 471 -633 477
rect -627 471 -624 477
rect -636 468 -624 471
rect -612 489 -600 498
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 477 -600 483
rect -612 471 -609 477
rect -603 471 -600 477
rect -612 468 -600 471
<< mvpdiff >>
rect -708 657 -696 660
rect -708 651 -705 657
rect -699 651 -696 657
rect -708 645 -696 651
rect -708 639 -705 645
rect -699 639 -696 645
rect -708 633 -696 639
rect -708 627 -705 633
rect -699 627 -696 633
rect -708 624 -696 627
rect -684 657 -672 660
rect -684 651 -681 657
rect -675 651 -672 657
rect -684 645 -672 651
rect -684 639 -681 645
rect -675 639 -672 645
rect -684 633 -672 639
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 624 -672 627
rect -660 657 -648 660
rect -660 651 -657 657
rect -651 651 -648 657
rect -660 645 -648 651
rect -660 639 -657 645
rect -651 639 -648 645
rect -660 633 -648 639
rect -660 627 -657 633
rect -651 627 -648 633
rect -660 624 -648 627
rect -636 657 -624 660
rect -636 651 -633 657
rect -627 651 -624 657
rect -636 645 -624 651
rect -636 639 -633 645
rect -627 639 -624 645
rect -636 633 -624 639
rect -636 627 -633 633
rect -627 627 -624 633
rect -636 624 -624 627
rect -612 657 -600 660
rect -612 651 -609 657
rect -603 651 -600 657
rect -612 645 -600 651
rect -612 639 -609 645
rect -603 639 -600 645
rect -612 633 -600 639
rect -612 627 -609 633
rect -603 627 -600 633
rect -612 624 -600 627
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -633 -81 -627 -75
rect -633 -93 -627 -87
rect -633 -105 -627 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
<< pdiffc >>
rect -705 483 -699 489
rect -705 471 -699 477
rect -681 483 -675 489
rect -681 471 -675 477
rect -657 483 -651 489
rect -657 471 -651 477
rect -633 483 -627 489
rect -633 471 -627 477
rect -609 483 -603 489
rect -609 471 -603 477
<< mvpdiffc >>
rect -705 651 -699 657
rect -705 639 -699 645
rect -705 627 -699 633
rect -681 651 -675 657
rect -681 639 -675 645
rect -681 627 -675 633
rect -657 651 -651 657
rect -657 639 -651 645
rect -657 627 -651 633
rect -633 651 -627 657
rect -633 639 -627 645
rect -633 627 -627 633
rect -609 651 -603 657
rect -609 639 -603 645
rect -609 627 -603 633
<< psubdiff >>
rect -720 705 -588 708
rect -720 699 -717 705
rect -711 699 -705 705
rect -699 699 -693 705
rect -687 699 -681 705
rect -675 699 -669 705
rect -663 699 -657 705
rect -651 699 -645 705
rect -639 699 -633 705
rect -627 699 -621 705
rect -615 699 -609 705
rect -603 699 -597 705
rect -591 699 -588 705
rect -720 696 -588 699
rect -720 561 -588 564
rect -720 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -657 561
rect -651 555 -645 561
rect -639 555 -633 561
rect -627 555 -621 561
rect -615 555 -609 561
rect -603 555 -597 561
rect -591 555 -588 561
rect -720 552 -588 555
rect -720 405 -588 408
rect -720 399 -717 405
rect -711 399 -705 405
rect -699 399 -693 405
rect -687 399 -681 405
rect -675 399 -669 405
rect -663 399 -657 405
rect -651 399 -645 405
rect -639 399 -633 405
rect -627 399 -621 405
rect -615 399 -609 405
rect -603 399 -597 405
rect -591 399 -588 405
rect -720 396 -588 399
rect -720 285 -588 288
rect -720 279 -717 285
rect -711 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -669 285
rect -663 279 -657 285
rect -651 279 -645 285
rect -639 279 -633 285
rect -627 279 -621 285
rect -615 279 -609 285
rect -603 279 -597 285
rect -591 279 -588 285
rect -720 276 -588 279
rect -720 237 -588 240
rect -720 231 -717 237
rect -711 231 -705 237
rect -699 231 -693 237
rect -687 231 -681 237
rect -675 231 -669 237
rect -663 231 -657 237
rect -651 231 -645 237
rect -639 231 -633 237
rect -627 231 -621 237
rect -615 231 -609 237
rect -603 231 -597 237
rect -591 231 -588 237
rect -720 228 -588 231
rect -720 189 -588 192
rect -720 183 -717 189
rect -711 183 -705 189
rect -699 183 -693 189
rect -687 183 -681 189
rect -675 183 -669 189
rect -663 183 -657 189
rect -651 183 -645 189
rect -639 183 -633 189
rect -627 183 -621 189
rect -615 183 -609 189
rect -603 183 -597 189
rect -591 183 -588 189
rect -720 180 -588 183
rect -720 141 -588 144
rect -720 135 -717 141
rect -711 135 -705 141
rect -699 135 -693 141
rect -687 135 -681 141
rect -675 135 -669 141
rect -663 135 -657 141
rect -651 135 -645 141
rect -639 135 -633 141
rect -627 135 -621 141
rect -615 135 -609 141
rect -603 135 -597 141
rect -591 135 -588 141
rect -720 132 -588 135
rect -720 93 -588 96
rect -720 87 -717 93
rect -711 87 -705 93
rect -699 87 -693 93
rect -687 87 -681 93
rect -675 87 -669 93
rect -663 87 -657 93
rect -651 87 -645 93
rect -639 87 -633 93
rect -627 87 -621 93
rect -615 87 -609 93
rect -603 87 -597 93
rect -591 87 -588 93
rect -720 84 -588 87
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< nsubdiff >>
rect -708 537 -600 540
rect -708 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -669 537
rect -663 531 -657 537
rect -651 531 -645 537
rect -639 531 -633 537
rect -627 531 -621 537
rect -615 531 -609 537
rect -603 531 -600 537
rect -708 528 -600 531
rect -708 429 -600 432
rect -708 423 -705 429
rect -699 423 -693 429
rect -687 423 -681 429
rect -675 423 -669 429
rect -663 423 -657 429
rect -651 423 -645 429
rect -639 423 -633 429
rect -627 423 -621 429
rect -615 423 -609 429
rect -603 423 -600 429
rect -708 420 -600 423
<< mvnsubdiff >>
rect -708 681 -600 684
rect -708 675 -705 681
rect -699 675 -693 681
rect -687 675 -681 681
rect -675 675 -669 681
rect -663 675 -657 681
rect -651 675 -645 681
rect -639 675 -633 681
rect -627 675 -621 681
rect -615 675 -609 681
rect -603 675 -600 681
rect -708 672 -600 675
rect -708 585 -600 588
rect -708 579 -705 585
rect -699 579 -693 585
rect -687 579 -681 585
rect -675 579 -669 585
rect -663 579 -657 585
rect -651 579 -645 585
rect -639 579 -633 585
rect -627 579 -621 585
rect -615 579 -609 585
rect -603 579 -600 585
rect -708 576 -600 579
<< psubdiffcont >>
rect -717 699 -711 705
rect -705 699 -699 705
rect -693 699 -687 705
rect -681 699 -675 705
rect -669 699 -663 705
rect -657 699 -651 705
rect -645 699 -639 705
rect -633 699 -627 705
rect -621 699 -615 705
rect -609 699 -603 705
rect -597 699 -591 705
rect -717 555 -711 561
rect -705 555 -699 561
rect -693 555 -687 561
rect -681 555 -675 561
rect -669 555 -663 561
rect -657 555 -651 561
rect -645 555 -639 561
rect -633 555 -627 561
rect -621 555 -615 561
rect -609 555 -603 561
rect -597 555 -591 561
rect -717 399 -711 405
rect -705 399 -699 405
rect -693 399 -687 405
rect -681 399 -675 405
rect -669 399 -663 405
rect -657 399 -651 405
rect -645 399 -639 405
rect -633 399 -627 405
rect -621 399 -615 405
rect -609 399 -603 405
rect -597 399 -591 405
rect -717 279 -711 285
rect -705 279 -699 285
rect -693 279 -687 285
rect -681 279 -675 285
rect -669 279 -663 285
rect -657 279 -651 285
rect -645 279 -639 285
rect -633 279 -627 285
rect -621 279 -615 285
rect -609 279 -603 285
rect -597 279 -591 285
rect -717 231 -711 237
rect -705 231 -699 237
rect -693 231 -687 237
rect -681 231 -675 237
rect -669 231 -663 237
rect -657 231 -651 237
rect -645 231 -639 237
rect -633 231 -627 237
rect -621 231 -615 237
rect -609 231 -603 237
rect -597 231 -591 237
rect -717 183 -711 189
rect -705 183 -699 189
rect -693 183 -687 189
rect -681 183 -675 189
rect -669 183 -663 189
rect -657 183 -651 189
rect -645 183 -639 189
rect -633 183 -627 189
rect -621 183 -615 189
rect -609 183 -603 189
rect -597 183 -591 189
rect -717 135 -711 141
rect -705 135 -699 141
rect -693 135 -687 141
rect -681 135 -675 141
rect -669 135 -663 141
rect -657 135 -651 141
rect -645 135 -639 141
rect -633 135 -627 141
rect -621 135 -615 141
rect -609 135 -603 141
rect -597 135 -591 141
rect -717 87 -711 93
rect -705 87 -699 93
rect -693 87 -687 93
rect -681 87 -675 93
rect -669 87 -663 93
rect -657 87 -651 93
rect -645 87 -639 93
rect -633 87 -627 93
rect -621 87 -615 93
rect -609 87 -603 93
rect -597 87 -591 93
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -657 -33 -651 -27
rect -645 -33 -639 -27
rect -633 -33 -627 -27
rect -621 -33 -615 -27
rect -609 -33 -603 -27
rect -597 -33 -591 -27
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
rect -657 -129 -651 -123
rect -645 -129 -639 -123
rect -633 -129 -627 -123
rect -621 -129 -615 -123
rect -609 -129 -603 -123
rect -597 -129 -591 -123
<< nsubdiffcont >>
rect -705 531 -699 537
rect -693 531 -687 537
rect -681 531 -675 537
rect -669 531 -663 537
rect -657 531 -651 537
rect -645 531 -639 537
rect -633 531 -627 537
rect -621 531 -615 537
rect -609 531 -603 537
rect -705 423 -699 429
rect -693 423 -687 429
rect -681 423 -675 429
rect -669 423 -663 429
rect -657 423 -651 429
rect -645 423 -639 429
rect -633 423 -627 429
rect -621 423 -615 429
rect -609 423 -603 429
<< mvnsubdiffcont >>
rect -705 675 -699 681
rect -693 675 -687 681
rect -681 675 -675 681
rect -669 675 -663 681
rect -657 675 -651 681
rect -645 675 -639 681
rect -633 675 -627 681
rect -621 675 -615 681
rect -609 675 -603 681
rect -705 579 -699 585
rect -693 579 -687 585
rect -681 579 -675 585
rect -669 579 -663 585
rect -657 579 -651 585
rect -645 579 -639 585
rect -633 579 -627 585
rect -621 579 -615 585
rect -609 579 -603 585
<< polysilicon >>
rect -696 660 -684 666
rect -672 660 -660 666
rect -648 660 -636 666
rect -624 660 -612 666
rect -696 612 -684 624
rect -672 612 -660 624
rect -648 612 -636 624
rect -624 612 -612 624
rect -696 609 -612 612
rect -696 603 -693 609
rect -687 603 -681 609
rect -675 603 -669 609
rect -663 603 -657 609
rect -651 603 -645 609
rect -639 603 -633 609
rect -627 603 -621 609
rect -615 603 -612 609
rect -696 600 -612 603
rect -696 498 -684 504
rect -672 498 -660 504
rect -648 498 -636 504
rect -624 498 -612 504
rect -696 456 -684 468
rect -672 456 -660 468
rect -696 453 -660 456
rect -696 447 -693 453
rect -687 447 -681 453
rect -675 447 -669 453
rect -663 447 -660 453
rect -696 444 -660 447
rect -648 456 -636 468
rect -624 456 -612 468
rect -648 453 -612 456
rect -648 447 -645 453
rect -639 447 -633 453
rect -627 447 -621 453
rect -615 447 -612 453
rect -648 444 -612 447
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -696 -72 -684 -60
rect -672 -72 -660 -60
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -648 -72 -636 -60
rect -624 -72 -612 -60
rect -696 -114 -684 -108
rect -672 -114 -660 -108
rect -648 -114 -636 -108
rect -624 -114 -612 -108
<< polycontact >>
rect -693 603 -687 609
rect -681 603 -675 609
rect -669 603 -663 609
rect -657 603 -651 609
rect -645 603 -639 609
rect -633 603 -627 609
rect -621 603 -615 609
rect -693 447 -687 453
rect -681 447 -675 453
rect -669 447 -663 453
rect -645 447 -639 453
rect -633 447 -627 453
rect -621 447 -615 453
rect -693 -57 -687 -51
rect -681 -57 -675 -51
rect -669 -57 -663 -51
rect -645 -57 -639 -51
rect -633 -57 -627 -51
rect -621 -57 -615 -51
<< metal1 >>
rect -720 705 -588 708
rect -720 699 -717 705
rect -711 699 -705 705
rect -699 699 -693 705
rect -687 699 -681 705
rect -675 699 -669 705
rect -663 699 -657 705
rect -651 699 -645 705
rect -639 699 -633 705
rect -627 699 -621 705
rect -615 699 -609 705
rect -603 699 -597 705
rect -591 699 -588 705
rect -720 696 -588 699
rect -720 681 -588 684
rect -720 675 -705 681
rect -699 675 -693 681
rect -687 675 -681 681
rect -675 675 -669 681
rect -663 675 -657 681
rect -651 675 -645 681
rect -639 675 -633 681
rect -627 675 -621 681
rect -615 675 -609 681
rect -603 675 -588 681
rect -720 672 -588 675
rect -708 657 -696 660
rect -708 651 -705 657
rect -699 651 -696 657
rect -708 645 -696 651
rect -708 639 -705 645
rect -699 639 -696 645
rect -708 633 -696 639
rect -708 627 -705 633
rect -699 627 -696 633
rect -708 624 -696 627
rect -684 657 -672 660
rect -684 651 -681 657
rect -675 651 -672 657
rect -684 645 -672 651
rect -684 639 -681 645
rect -675 639 -672 645
rect -684 633 -672 639
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 624 -672 627
rect -660 657 -648 660
rect -660 651 -657 657
rect -651 651 -648 657
rect -660 645 -648 651
rect -660 639 -657 645
rect -651 639 -648 645
rect -660 633 -648 639
rect -660 627 -657 633
rect -651 627 -648 633
rect -660 624 -648 627
rect -636 657 -624 660
rect -636 651 -633 657
rect -627 651 -624 657
rect -636 645 -624 651
rect -636 639 -633 645
rect -627 639 -624 645
rect -636 633 -624 639
rect -636 627 -633 633
rect -627 627 -624 633
rect -636 624 -624 627
rect -612 657 -600 660
rect -612 651 -609 657
rect -603 651 -600 657
rect -612 645 -600 651
rect -612 639 -609 645
rect -603 639 -600 645
rect -612 633 -600 639
rect -612 627 -609 633
rect -603 627 -600 633
rect -612 624 -600 627
rect -696 609 -612 612
rect -696 603 -693 609
rect -687 603 -681 609
rect -675 603 -669 609
rect -663 603 -657 609
rect -651 603 -645 609
rect -639 603 -633 609
rect -627 603 -621 609
rect -615 603 -612 609
rect -696 600 -612 603
rect -720 585 -588 588
rect -720 579 -705 585
rect -699 579 -693 585
rect -687 579 -681 585
rect -675 579 -669 585
rect -663 579 -657 585
rect -651 579 -645 585
rect -639 579 -633 585
rect -627 579 -621 585
rect -615 579 -609 585
rect -603 579 -588 585
rect -720 576 -588 579
rect -720 561 -588 564
rect -720 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -657 561
rect -651 555 -645 561
rect -639 555 -633 561
rect -627 555 -621 561
rect -615 555 -609 561
rect -603 555 -597 561
rect -591 555 -588 561
rect -720 552 -588 555
rect -720 537 -588 540
rect -720 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -669 537
rect -663 531 -657 537
rect -651 531 -645 537
rect -639 531 -633 537
rect -627 531 -621 537
rect -615 531 -609 537
rect -603 531 -588 537
rect -720 528 -588 531
rect -708 513 -600 516
rect -708 507 -705 513
rect -699 507 -657 513
rect -651 507 -609 513
rect -603 507 -600 513
rect -708 504 -600 507
rect -708 501 -696 504
rect -708 495 -705 501
rect -699 495 -696 501
rect -660 501 -648 504
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 477 -696 483
rect -708 471 -705 477
rect -699 471 -696 477
rect -708 468 -696 471
rect -684 489 -672 498
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 477 -672 483
rect -684 471 -681 477
rect -675 471 -672 477
rect -684 468 -672 471
rect -660 495 -657 501
rect -651 495 -648 501
rect -612 501 -600 504
rect -660 489 -648 495
rect -660 483 -657 489
rect -651 483 -648 489
rect -660 477 -648 483
rect -660 471 -657 477
rect -651 471 -648 477
rect -660 468 -648 471
rect -636 489 -624 498
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 477 -624 483
rect -636 471 -633 477
rect -627 471 -624 477
rect -636 468 -624 471
rect -612 495 -609 501
rect -603 495 -600 501
rect -612 489 -600 495
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 477 -600 483
rect -612 471 -609 477
rect -603 471 -600 477
rect -612 468 -600 471
rect -696 453 -660 456
rect -696 447 -693 453
rect -687 447 -681 453
rect -675 447 -669 453
rect -663 447 -660 453
rect -696 444 -660 447
rect -648 453 -612 456
rect -648 447 -645 453
rect -639 447 -633 453
rect -627 447 -621 453
rect -615 447 -612 453
rect -648 444 -612 447
rect -720 429 -588 432
rect -720 423 -705 429
rect -699 423 -693 429
rect -687 423 -681 429
rect -675 423 -669 429
rect -663 423 -657 429
rect -651 423 -645 429
rect -639 423 -633 429
rect -627 423 -621 429
rect -615 423 -609 429
rect -603 423 -588 429
rect -720 420 -588 423
rect -720 405 -588 408
rect -720 399 -717 405
rect -711 399 -705 405
rect -699 399 -693 405
rect -687 399 -681 405
rect -675 399 -669 405
rect -663 399 -657 405
rect -651 399 -645 405
rect -639 399 -633 405
rect -627 399 -621 405
rect -615 399 -609 405
rect -603 399 -597 405
rect -591 399 -588 405
rect -720 396 -588 399
rect -720 285 -588 288
rect -720 279 -717 285
rect -711 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -669 285
rect -663 279 -657 285
rect -651 279 -645 285
rect -639 279 -633 285
rect -627 279 -621 285
rect -615 279 -609 285
rect -603 279 -597 285
rect -591 279 -588 285
rect -720 276 -588 279
rect -720 237 -588 240
rect -720 231 -717 237
rect -711 231 -705 237
rect -699 231 -693 237
rect -687 231 -681 237
rect -675 231 -669 237
rect -663 231 -657 237
rect -651 231 -645 237
rect -639 231 -633 237
rect -627 231 -621 237
rect -615 231 -609 237
rect -603 231 -597 237
rect -591 231 -588 237
rect -720 228 -588 231
rect -720 189 -588 192
rect -720 183 -717 189
rect -711 183 -705 189
rect -699 183 -693 189
rect -687 183 -681 189
rect -675 183 -669 189
rect -663 183 -657 189
rect -651 183 -645 189
rect -639 183 -633 189
rect -627 183 -621 189
rect -615 183 -609 189
rect -603 183 -597 189
rect -591 183 -588 189
rect -720 180 -588 183
rect -720 141 -588 144
rect -720 135 -717 141
rect -711 135 -705 141
rect -699 135 -693 141
rect -687 135 -681 141
rect -675 135 -669 141
rect -663 135 -657 141
rect -651 135 -645 141
rect -639 135 -633 141
rect -627 135 -621 141
rect -615 135 -609 141
rect -603 135 -597 141
rect -591 135 -588 141
rect -720 132 -588 135
rect -720 93 -588 96
rect -720 87 -717 93
rect -711 87 -705 93
rect -699 87 -693 93
rect -687 87 -681 93
rect -675 87 -669 93
rect -663 87 -657 93
rect -651 87 -645 93
rect -639 87 -633 93
rect -627 87 -621 93
rect -615 87 -609 93
rect -603 87 -597 93
rect -591 87 -588 93
rect -720 84 -588 87
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< via1 >>
rect -705 675 -699 681
rect -657 675 -651 681
rect -609 675 -603 681
rect -705 651 -699 657
rect -705 639 -699 645
rect -705 627 -699 633
rect -681 651 -675 657
rect -681 639 -675 645
rect -681 627 -675 633
rect -657 651 -651 657
rect -657 639 -651 645
rect -657 627 -651 633
rect -633 651 -627 657
rect -633 639 -627 645
rect -633 627 -627 633
rect -609 651 -603 657
rect -609 639 -603 645
rect -609 627 -603 633
rect -657 603 -651 609
rect -705 507 -699 513
rect -657 507 -651 513
rect -609 507 -603 513
rect -705 495 -699 501
rect -705 483 -699 489
rect -705 471 -699 477
rect -681 483 -675 489
rect -681 471 -675 477
rect -657 495 -651 501
rect -633 483 -627 489
rect -633 471 -627 477
rect -609 495 -603 501
rect -609 483 -603 489
rect -609 471 -603 477
rect -681 447 -675 453
rect -633 447 -627 453
rect -705 423 -699 429
rect -609 423 -603 429
rect -705 399 -699 405
rect -609 399 -603 405
rect -705 279 -699 285
rect -609 279 -603 285
rect -705 231 -699 237
rect -609 231 -603 237
rect -705 183 -699 189
rect -609 183 -603 189
rect -705 135 -699 141
rect -609 135 -603 141
rect -705 87 -699 93
rect -609 87 -603 93
rect -705 -33 -699 -27
rect -609 -33 -603 -27
rect -681 -57 -675 -51
rect -633 -57 -627 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal2 >>
rect -708 681 -696 684
rect -708 675 -705 681
rect -699 675 -696 681
rect -708 657 -696 675
rect -660 681 -648 684
rect -660 675 -657 681
rect -651 675 -648 681
rect -708 651 -705 657
rect -699 651 -696 657
rect -708 645 -696 651
rect -708 639 -705 645
rect -699 639 -696 645
rect -708 633 -696 639
rect -708 627 -705 633
rect -699 627 -696 633
rect -708 624 -696 627
rect -684 657 -672 660
rect -684 651 -681 657
rect -675 651 -672 657
rect -684 645 -672 651
rect -684 639 -681 645
rect -675 639 -672 645
rect -684 633 -672 639
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 585 -672 627
rect -660 657 -648 675
rect -612 681 -600 684
rect -612 675 -609 681
rect -603 675 -600 681
rect -660 651 -657 657
rect -651 651 -648 657
rect -660 645 -648 651
rect -660 639 -657 645
rect -651 639 -648 645
rect -660 633 -648 639
rect -660 627 -657 633
rect -651 627 -648 633
rect -660 624 -648 627
rect -636 657 -624 660
rect -636 651 -633 657
rect -627 651 -624 657
rect -636 645 -624 651
rect -636 639 -633 645
rect -627 639 -624 645
rect -636 633 -624 639
rect -636 627 -633 633
rect -627 627 -624 633
rect -660 609 -648 612
rect -660 603 -657 609
rect -651 603 -648 609
rect -660 600 -648 603
rect -684 579 -681 585
rect -675 579 -672 585
rect -708 537 -696 540
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 513 -696 531
rect -684 537 -672 579
rect -636 585 -624 627
rect -612 657 -600 675
rect -612 651 -609 657
rect -603 651 -600 657
rect -612 645 -600 651
rect -612 639 -609 645
rect -603 639 -600 645
rect -612 633 -600 639
rect -612 627 -609 633
rect -603 627 -600 633
rect -612 624 -600 627
rect -636 579 -633 585
rect -627 579 -624 585
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 528 -672 531
rect -660 537 -648 540
rect -660 531 -657 537
rect -651 531 -648 537
rect -708 507 -705 513
rect -699 507 -696 513
rect -708 501 -696 507
rect -708 495 -705 501
rect -699 495 -696 501
rect -660 513 -648 531
rect -636 537 -624 579
rect -636 531 -633 537
rect -627 531 -624 537
rect -636 528 -624 531
rect -612 537 -600 540
rect -612 531 -609 537
rect -603 531 -600 537
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 501 -648 507
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 477 -696 483
rect -708 471 -705 477
rect -699 471 -696 477
rect -708 468 -696 471
rect -684 489 -672 498
rect -660 495 -657 501
rect -651 495 -648 501
rect -612 513 -600 531
rect -612 507 -609 513
rect -603 507 -600 513
rect -612 501 -600 507
rect -660 492 -648 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -636 489 -624 498
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 480 -624 483
rect -684 477 -624 480
rect -684 471 -681 477
rect -675 471 -633 477
rect -627 471 -624 477
rect -684 468 -624 471
rect -612 495 -609 501
rect -603 495 -600 501
rect -612 489 -600 495
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 477 -600 483
rect -612 471 -609 477
rect -603 471 -600 477
rect -612 468 -600 471
rect -684 453 -672 456
rect -684 447 -681 453
rect -675 447 -672 453
rect -684 444 -672 447
rect -708 429 -696 432
rect -708 423 -705 429
rect -699 423 -696 429
rect -708 420 -696 423
rect -708 405 -696 408
rect -708 399 -705 405
rect -699 399 -696 405
rect -708 285 -696 399
rect -708 279 -705 285
rect -699 279 -696 285
rect -708 237 -696 279
rect -708 231 -705 237
rect -699 231 -696 237
rect -708 189 -696 231
rect -708 183 -705 189
rect -699 183 -696 189
rect -708 141 -696 183
rect -708 135 -705 141
rect -699 135 -696 141
rect -708 93 -696 135
rect -708 87 -705 93
rect -699 87 -696 93
rect -708 -27 -696 87
rect -708 -33 -705 -27
rect -699 -33 -696 -27
rect -708 -75 -696 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -123 -696 -105
rect -660 -75 -648 468
rect -636 453 -624 456
rect -636 447 -633 453
rect -627 447 -624 453
rect -636 444 -624 447
rect -612 429 -600 432
rect -612 423 -609 429
rect -603 423 -600 429
rect -612 420 -600 423
rect -612 405 -600 408
rect -612 399 -609 405
rect -603 399 -600 405
rect -612 285 -600 399
rect -612 279 -609 285
rect -603 279 -600 285
rect -612 237 -600 279
rect -612 231 -609 237
rect -603 231 -600 237
rect -612 189 -600 231
rect -612 183 -609 189
rect -603 183 -600 189
rect -612 141 -600 183
rect -612 135 -609 141
rect -603 135 -600 141
rect -612 93 -600 135
rect -612 87 -609 93
rect -603 87 -600 93
rect -612 -27 -600 87
rect -612 -33 -609 -27
rect -603 -33 -600 -27
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -612 -75 -600 -33
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -708 -129 -705 -123
rect -699 -129 -696 -123
rect -708 -132 -696 -129
rect -612 -123 -600 -105
rect -612 -129 -609 -123
rect -603 -129 -600 -123
rect -612 -132 -600 -129
<< via2 >>
rect -705 675 -699 681
rect -657 675 -651 681
rect -705 651 -699 657
rect -705 639 -699 645
rect -705 627 -699 633
rect -609 675 -603 681
rect -657 651 -651 657
rect -657 639 -651 645
rect -657 627 -651 633
rect -657 603 -651 609
rect -681 579 -675 585
rect -705 531 -699 537
rect -609 651 -603 657
rect -609 639 -603 645
rect -609 627 -603 633
rect -633 579 -627 585
rect -681 531 -675 537
rect -657 531 -651 537
rect -633 531 -627 537
rect -609 531 -603 537
rect -681 447 -675 453
rect -705 423 -699 429
rect -705 399 -699 405
rect -705 279 -699 285
rect -705 231 -699 237
rect -705 183 -699 189
rect -705 135 -699 141
rect -705 87 -699 93
rect -705 -33 -699 -27
rect -681 -57 -675 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -633 447 -627 453
rect -609 423 -603 429
rect -609 399 -603 405
rect -609 279 -603 285
rect -609 231 -603 237
rect -609 183 -603 189
rect -609 135 -603 141
rect -609 87 -603 93
rect -609 -33 -603 -27
rect -633 -57 -627 -51
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal3 >>
rect -720 681 -588 684
rect -720 675 -705 681
rect -699 675 -657 681
rect -651 675 -609 681
rect -603 675 -588 681
rect -720 657 -588 675
rect -720 651 -705 657
rect -699 651 -657 657
rect -651 651 -609 657
rect -603 651 -588 657
rect -720 645 -588 651
rect -720 639 -705 645
rect -699 639 -657 645
rect -651 639 -609 645
rect -603 639 -588 645
rect -720 633 -588 639
rect -720 627 -705 633
rect -699 627 -657 633
rect -651 627 -609 633
rect -603 627 -588 633
rect -720 624 -588 627
rect -660 609 -648 612
rect -660 603 -657 609
rect -651 603 -648 609
rect -660 600 -648 603
rect -720 585 -588 588
rect -720 579 -681 585
rect -675 579 -633 585
rect -627 579 -588 585
rect -720 570 -588 579
rect -720 561 -588 564
rect -720 555 -657 561
rect -651 555 -588 561
rect -720 552 -588 555
rect -720 537 -588 546
rect -720 531 -705 537
rect -699 531 -681 537
rect -675 531 -657 537
rect -651 531 -633 537
rect -627 531 -609 537
rect -603 531 -588 537
rect -720 528 -588 531
rect -684 453 -672 456
rect -684 447 -681 453
rect -675 447 -672 453
rect -684 444 -672 447
rect -636 453 -624 456
rect -636 447 -633 453
rect -627 447 -624 453
rect -636 444 -624 447
rect -720 429 -588 432
rect -720 423 -705 429
rect -699 423 -609 429
rect -603 423 -588 429
rect -720 420 -588 423
rect -720 405 -588 408
rect -720 399 -705 405
rect -699 399 -609 405
rect -603 399 -588 405
rect -720 396 -588 399
rect -720 354 -588 384
rect -720 336 -588 348
rect -720 300 -588 330
rect -720 285 -588 288
rect -720 279 -705 285
rect -699 279 -609 285
rect -603 279 -588 285
rect -720 276 -588 279
rect -720 252 -588 264
rect -720 237 -588 240
rect -720 231 -705 237
rect -699 231 -609 237
rect -603 231 -588 237
rect -720 228 -588 231
rect -720 204 -588 216
rect -720 189 -588 192
rect -720 183 -705 189
rect -699 183 -609 189
rect -603 183 -588 189
rect -720 180 -588 183
rect -720 156 -588 168
rect -720 141 -588 144
rect -720 135 -705 141
rect -699 135 -609 141
rect -603 135 -588 141
rect -720 132 -588 135
rect -720 108 -588 120
rect -720 93 -588 96
rect -720 87 -705 93
rect -699 87 -609 93
rect -603 87 -588 93
rect -720 84 -588 87
rect -720 42 -588 72
rect -720 24 -588 36
rect -720 -12 -588 18
rect -720 -27 -588 -24
rect -720 -33 -705 -27
rect -699 -33 -609 -27
rect -603 -33 -588 -27
rect -720 -36 -588 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -720 -75 -588 -72
rect -720 -81 -705 -75
rect -699 -81 -609 -75
rect -603 -81 -588 -75
rect -720 -87 -588 -81
rect -720 -93 -705 -87
rect -699 -93 -609 -87
rect -603 -93 -588 -87
rect -720 -99 -588 -93
rect -720 -105 -705 -99
rect -699 -105 -609 -99
rect -603 -105 -588 -99
rect -720 -123 -588 -105
rect -720 -129 -705 -123
rect -699 -129 -609 -123
rect -603 -129 -588 -123
rect -720 -132 -588 -129
<< via3 >>
rect -657 603 -651 609
rect -681 579 -675 585
rect -633 579 -627 585
rect -657 555 -651 561
rect -705 531 -699 537
rect -681 531 -675 537
rect -633 531 -627 537
rect -609 531 -603 537
rect -681 447 -675 453
rect -633 447 -627 453
rect -681 -57 -675 -51
rect -633 -57 -627 -51
<< metal4 >>
rect -660 609 -648 612
rect -660 603 -657 609
rect -651 603 -648 609
rect -684 585 -672 588
rect -684 579 -681 585
rect -675 579 -672 585
rect -708 537 -696 540
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 528 -696 531
rect -684 537 -672 579
rect -660 561 -648 603
rect -660 555 -657 561
rect -651 555 -648 561
rect -660 552 -648 555
rect -636 585 -624 588
rect -636 579 -633 585
rect -627 579 -624 585
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 528 -672 531
rect -636 537 -624 579
rect -636 531 -633 537
rect -627 531 -624 537
rect -636 528 -624 531
rect -612 537 -600 540
rect -612 531 -609 537
rect -603 531 -600 537
rect -612 528 -600 531
rect -684 453 -672 456
rect -684 447 -681 453
rect -675 447 -672 453
rect -684 432 -672 447
rect -708 420 -672 432
rect -684 -51 -672 420
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 453 -624 456
rect -636 447 -633 453
rect -627 447 -624 453
rect -636 432 -624 447
rect -636 420 -600 432
rect -636 -51 -624 420
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
<< labels >>
rlabel metal4 -684 -12 -672 240 0 inl
port 1 nsew
rlabel metal4 -636 -12 -624 240 0 inr
port 2 nsew
rlabel metal2 -660 -12 -648 240 0 out
port 3 nsew
rlabel metal3 -720 -132 -588 -72 0 gnd
port 14 nsew
rlabel metal1 -684 -108 -672 -72 0 dl
rlabel metal1 -636 -108 -624 -72 0 dr
rlabel metal3 -720 -12 -588 0 0 om
port 15 nsew
rlabel metal3 -720 24 -588 36 0 xp
port 13 nsew
rlabel metal3 -720 108 -588 120 0 ip
port 11 nsew
rlabel metal3 -720 60 -588 72 0 om
port 15 nsew
rlabel metal3 -720 252 -588 264 0 im
port 10 nsew
rlabel metal3 -720 336 -588 348 0 xm
port 9 nsew
rlabel metal3 -720 624 -588 684 0 vdd
port 4 nsew
rlabel metal3 -720 552 -708 564 0 gp
port 5 nsew
rlabel metal3 -720 420 -708 432 0 bp
port 6 nsew
rlabel metal3 -720 576 -708 588 0 vreg
port 7 nsew
rlabel metal3 -720 372 -588 384 0 op
port 8 nsew
rlabel metal1 -708 552 -696 564 0 gnd
rlabel metal1 -708 696 -696 708 0 gnd
rlabel metal3 -720 300 -588 312 0 op
port 8 nsew
rlabel metal3 -720 204 -588 216 0 x
port 16 nsew
rlabel metal3 -720 156 -588 168 0 y
port 17 nsew
<< end >>
