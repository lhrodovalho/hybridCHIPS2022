magic
tech gf180mcuC
magscale 1 5
timestamp 1665299795
<< metal1 >>
rect -5040 1440 -4980 1500
rect 2760 1440 2820 1500
<< metal2 >>
rect -4440 1254 -4380 1260
rect -4440 966 -4424 1254
rect -4396 966 -4380 1254
rect -4440 960 -4380 966
rect -1440 1254 -1380 1260
rect -1440 966 -1424 1254
rect -1396 966 -1380 1254
rect -1440 960 -1380 966
rect -840 1254 -780 1260
rect -840 966 -824 1254
rect -796 966 -780 1254
rect -840 960 -780 966
rect 2160 1254 2220 1260
rect 2160 966 2176 1254
rect 2204 966 2220 1254
rect 2160 960 2220 966
rect -3240 524 -3180 540
rect -3240 496 -3224 524
rect -3196 496 -3180 524
rect -3240 480 -3180 496
rect -2640 524 -2580 540
rect -2640 496 -2624 524
rect -2596 496 -2580 524
rect -2640 480 -2580 496
rect 360 524 420 540
rect 360 496 376 524
rect 404 496 420 524
rect 360 480 420 496
rect 960 524 1020 540
rect 960 496 976 524
rect 1004 496 1020 524
rect 960 480 1020 496
rect -3840 54 -3780 60
rect -3840 -234 -3824 54
rect -3796 -234 -3780 54
rect -3840 -240 -3780 -234
rect -2040 54 -1980 60
rect -2040 -234 -2024 54
rect -1996 -234 -1980 54
rect -2040 -240 -1980 -234
rect -240 54 -180 60
rect -240 -234 -224 54
rect -196 -234 -180 54
rect -240 -240 -180 -234
rect 1560 54 1620 60
rect 1560 -234 1576 54
rect 1604 -234 1620 54
rect 1560 -240 1620 -234
<< via2 >>
rect -4424 966 -4396 1254
rect -1424 966 -1396 1254
rect -824 966 -796 1254
rect 2176 966 2204 1254
rect -3224 496 -3196 524
rect -2624 496 -2596 524
rect 376 496 404 524
rect 976 496 1004 524
rect -3824 -234 -3796 54
rect -2024 -234 -1996 54
rect -224 -234 -196 54
rect 1576 -234 1604 54
<< metal3 >>
rect -5220 2460 -5160 2760
rect -5220 2190 -5160 2280
rect -5220 2100 -5160 2160
rect -5220 1440 2940 1500
rect -5220 960 -5160 1260
rect -4440 1254 -4380 1260
rect -4440 966 -4424 1254
rect -4396 966 -4380 1254
rect -4440 960 -4380 966
rect -1440 1254 -1380 1260
rect -1440 966 -1424 1254
rect -1396 966 -1380 1254
rect -1440 960 -1380 966
rect -840 1254 -780 1260
rect -840 966 -824 1254
rect -796 966 -780 1254
rect -840 960 -780 966
rect 2160 1254 2220 1260
rect 2160 966 2176 1254
rect 2204 966 2220 1254
rect 2160 960 2220 966
rect -5220 720 -5160 780
rect -4560 764 -4500 780
rect -4560 736 -4544 764
rect -4516 736 -4500 764
rect -4560 720 -4500 736
rect -2520 764 -2460 780
rect -2520 736 -2504 764
rect -2476 736 -2460 764
rect -2520 720 -2460 736
rect -1320 764 -1260 780
rect -1320 736 -1304 764
rect -1276 736 -1260 764
rect -1320 720 -1260 736
rect -960 764 -900 780
rect -960 736 -944 764
rect -916 736 -900 764
rect -960 720 -900 736
rect 240 764 300 780
rect 240 736 256 764
rect 284 736 300 764
rect 240 720 300 736
rect 2280 764 2340 780
rect 2280 736 2296 764
rect 2324 736 2340 764
rect 2280 720 2340 736
rect -5220 480 -5160 540
rect -4320 524 -4260 540
rect -4320 496 -4304 524
rect -4276 496 -4260 524
rect -4320 480 -4260 496
rect -3960 524 -3900 540
rect -3960 496 -3944 524
rect -3916 496 -3900 524
rect -3960 480 -3900 496
rect -3240 524 -3180 540
rect -3240 496 -3224 524
rect -3196 496 -3180 524
rect -3240 480 -3180 496
rect -3120 524 -3060 540
rect -3120 496 -3104 524
rect -3076 496 -3060 524
rect -3120 480 -3060 496
rect -2760 524 -2700 540
rect -2760 496 -2744 524
rect -2716 496 -2700 524
rect -2760 480 -2700 496
rect -2640 524 -2580 540
rect -2640 496 -2624 524
rect -2596 496 -2580 524
rect -2640 480 -2580 496
rect -1920 524 -1860 540
rect -1920 496 -1904 524
rect -1876 496 -1860 524
rect -1920 480 -1860 496
rect -1560 524 -1500 540
rect -1560 496 -1544 524
rect -1516 496 -1500 524
rect -1560 480 -1500 496
rect -720 524 -660 540
rect -720 496 -704 524
rect -676 496 -660 524
rect -720 480 -660 496
rect -360 524 -300 540
rect -360 496 -344 524
rect -316 496 -300 524
rect -360 480 -300 496
rect 360 524 420 540
rect 360 496 376 524
rect 404 496 420 524
rect 360 480 420 496
rect 480 524 540 540
rect 480 496 496 524
rect 524 496 540 524
rect 480 480 540 496
rect 840 524 900 540
rect 840 496 856 524
rect 884 496 900 524
rect 840 480 900 496
rect 960 524 1020 540
rect 960 496 976 524
rect 1004 496 1020 524
rect 960 480 1020 496
rect 1680 524 1740 540
rect 1680 496 1696 524
rect 1724 496 1740 524
rect 1680 480 1740 496
rect 2040 524 2100 540
rect 2040 496 2056 524
rect 2084 496 2100 524
rect 2040 480 2100 496
rect -5220 240 -5160 300
rect -3720 284 -3660 300
rect -3720 256 -3704 284
rect -3676 256 -3660 284
rect -3720 240 -3660 256
rect -3360 284 -3300 300
rect -3360 256 -3344 284
rect -3316 256 -3300 284
rect -3360 240 -3300 256
rect -2160 284 -2100 300
rect -2160 256 -2144 284
rect -2116 256 -2100 284
rect -2160 240 -2100 256
rect -120 284 -60 300
rect -120 256 -104 284
rect -76 256 -60 284
rect -120 240 -60 256
rect 1080 284 1140 300
rect 1080 256 1096 284
rect 1124 256 1140 284
rect 1080 240 1140 256
rect 1440 284 1500 300
rect 1440 256 1456 284
rect 1484 256 1500 284
rect 1440 240 1500 256
rect -5220 -240 -5160 60
rect -3840 54 -3780 60
rect -3840 -234 -3824 54
rect -3796 -234 -3780 54
rect -3840 -240 -3780 -234
rect -2040 54 -1980 60
rect -2040 -234 -2024 54
rect -1996 -234 -1980 54
rect -2040 -240 -1980 -234
rect -240 54 -180 60
rect -240 -234 -224 54
rect -196 -234 -180 54
rect -240 -240 -180 -234
rect 1560 54 1620 60
rect 1560 -234 1576 54
rect 1604 -234 1620 54
rect 1560 -240 1620 -234
rect -5220 -840 -5160 -540
<< via3 >>
rect -4544 736 -4516 764
rect -2504 736 -2476 764
rect -1304 736 -1276 764
rect -944 736 -916 764
rect 256 736 284 764
rect 2296 736 2324 764
rect -4304 496 -4276 524
rect -3944 496 -3916 524
rect -3104 496 -3076 524
rect -2744 496 -2716 524
rect -1904 496 -1876 524
rect -1544 496 -1516 524
rect -704 496 -676 524
rect -344 496 -316 524
rect 496 496 524 524
rect 856 496 884 524
rect 1696 496 1724 524
rect 2056 496 2084 524
rect -3704 256 -3676 284
rect -3344 256 -3316 284
rect -2144 256 -2116 284
rect -104 256 -76 284
rect 1096 256 1124 284
rect 1456 256 1484 284
<< metal4 >>
rect -4560 764 -4500 780
rect -4560 736 -4544 764
rect -4516 736 -4500 764
rect -4560 720 -4500 736
rect -2520 764 -2460 780
rect -2520 736 -2504 764
rect -2476 736 -2460 764
rect -2520 720 -2460 736
rect -1320 764 -1260 780
rect -1320 736 -1304 764
rect -1276 736 -1260 764
rect -1320 720 -1260 736
rect -960 764 -900 780
rect -960 736 -944 764
rect -916 736 -900 764
rect -960 720 -900 736
rect 240 764 300 780
rect 240 736 256 764
rect 284 736 300 764
rect 240 720 300 736
rect 2280 764 2340 780
rect 2280 736 2296 764
rect 2324 736 2340 764
rect 2280 720 2340 736
rect -4320 524 -4260 540
rect -4320 496 -4304 524
rect -4276 496 -4260 524
rect -4320 480 -4260 496
rect -3960 524 -3900 540
rect -3960 496 -3944 524
rect -3916 496 -3900 524
rect -3960 480 -3900 496
rect -3120 524 -3060 540
rect -3120 496 -3104 524
rect -3076 496 -3060 524
rect -3120 480 -3060 496
rect -2760 524 -2700 540
rect -2760 496 -2744 524
rect -2716 496 -2700 524
rect -2760 480 -2700 496
rect -1920 524 -1860 540
rect -1920 496 -1904 524
rect -1876 496 -1860 524
rect -1920 480 -1860 496
rect -1560 524 -1500 540
rect -1560 496 -1544 524
rect -1516 496 -1500 524
rect -1560 480 -1500 496
rect -720 524 -660 540
rect -720 496 -704 524
rect -676 496 -660 524
rect -720 480 -660 496
rect -360 524 -300 540
rect -360 496 -344 524
rect -316 496 -300 524
rect -360 480 -300 496
rect 480 524 540 540
rect 480 496 496 524
rect 524 496 540 524
rect 480 480 540 496
rect 840 524 900 540
rect 840 496 856 524
rect 884 496 900 524
rect 840 480 900 496
rect 1680 524 1740 540
rect 1680 496 1696 524
rect 1724 496 1740 524
rect 1680 480 1740 496
rect 2040 524 2100 540
rect 2040 496 2056 524
rect 2084 496 2100 524
rect 2040 480 2100 496
rect -3720 284 -3660 300
rect -3720 256 -3704 284
rect -3676 256 -3660 284
rect -3720 240 -3660 256
rect -3360 284 -3300 300
rect -3360 256 -3344 284
rect -3316 256 -3300 284
rect -3360 240 -3300 256
rect -2160 284 -2100 300
rect -2160 256 -2144 284
rect -2116 256 -2100 284
rect -2160 240 -2100 256
rect -120 284 -60 300
rect -120 256 -104 284
rect -76 256 -60 284
rect -120 240 -60 256
rect 1080 284 1140 300
rect 1080 256 1096 284
rect 1124 256 1140 284
rect 1080 240 1140 256
rect 1440 284 1500 300
rect 1440 256 1456 284
rect 1484 256 1500 284
rect 1440 240 1500 256
use barth_cell#0  barth_cell_0
timestamp 1665184495
transform -1 0 -1080 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_1
timestamp 1665184495
transform -1 0 -1680 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_2
timestamp 1665184495
transform -1 0 -2280 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_3
timestamp 1665184495
transform -1 0 -2880 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_4
timestamp 1665184495
transform -1 0 -3480 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_5
timestamp 1665184495
transform -1 0 -4080 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_6
timestamp 1665184495
transform 1 0 1860 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_7
timestamp 1665184495
transform 1 0 1260 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_8
timestamp 1665184495
transform 1 0 660 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_9
timestamp 1665184495
transform 1 0 60 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_10
timestamp 1665184495
transform 1 0 -540 0 1 -180
box -3600 -660 -2940 3060
use barth_cell#0  barth_cell_11
timestamp 1665184495
transform 1 0 -1140 0 1 -180
box -3600 -660 -2940 3060
use barth_edge#0  barth_edge_0
timestamp 1665184495
transform -1 0 -840 0 1 -180
box -3780 -660 -3300 3060
use barth_edge#0  barth_edge_1
timestamp 1665184495
transform 1 0 -1380 0 1 -180
box -3780 -660 -3300 3060
<< labels >>
rlabel metal3 s -5190 510 -5190 510 4 x
rlabel metal3 s -5220 240 -5160 300 4 ip
port 1 nsew
rlabel metal3 s -5220 720 -5160 780 4 im
port 2 nsew
rlabel metal3 s -5220 960 -5160 1260 4 op
port 3 nsew
rlabel metal3 s -5220 -240 -5160 60 4 om
port 4 nsew
rlabel metal3 s -5220 2460 -5160 2760 4 vdd
port 5 nsew
rlabel metal3 s -5220 2100 -5160 2160 4 gp
port 6 nsew
rlabel metal3 s -5220 1440 -5160 1500 4 bp
port 7 nsew
rlabel metal3 s -5220 2220 -5160 2280 4 vreg
port 8 nsew
rlabel metal3 s -5220 -840 -5160 -540 4 gnd
port 9 nsew
<< end >>
