magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7200 4740 -5880 5940
rect -7200 3180 -5880 4500
<< nmos >>
rect -6960 -1080 -6840 -720
rect -6720 -1080 -6600 -720
rect -6480 -1080 -6360 -720
rect -6240 -1080 -6120 -720
<< pmos >>
rect -6960 3720 -6840 4020
rect -6720 3720 -6600 4020
rect -6480 3720 -6360 4020
rect -6240 3720 -6120 4020
<< mvpmos >>
rect -6960 5280 -6840 5640
rect -6720 5280 -6600 5640
rect -6480 5280 -6360 5640
rect -6240 5280 -6120 5640
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -757 -6480 -720
rect -6600 -803 -6563 -757
rect -6517 -803 -6480 -757
rect -6600 -877 -6480 -803
rect -6600 -923 -6563 -877
rect -6517 -923 -6480 -877
rect -6600 -997 -6480 -923
rect -6600 -1043 -6563 -997
rect -6517 -1043 -6480 -997
rect -6600 -1080 -6480 -1043
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -757 -6000 -720
rect -6120 -803 -6083 -757
rect -6037 -803 -6000 -757
rect -6120 -877 -6000 -803
rect -6120 -923 -6083 -877
rect -6037 -923 -6000 -877
rect -6120 -997 -6000 -923
rect -6120 -1043 -6083 -997
rect -6037 -1043 -6000 -997
rect -6120 -1080 -6000 -1043
<< pdiff >>
rect -7080 3923 -6960 4020
rect -7080 3877 -7043 3923
rect -6997 3877 -6960 3923
rect -7080 3803 -6960 3877
rect -7080 3757 -7043 3803
rect -6997 3757 -6960 3803
rect -7080 3720 -6960 3757
rect -6840 3923 -6720 4020
rect -6840 3877 -6803 3923
rect -6757 3877 -6720 3923
rect -6840 3803 -6720 3877
rect -6840 3757 -6803 3803
rect -6757 3757 -6720 3803
rect -6840 3720 -6720 3757
rect -6600 3923 -6480 4020
rect -6600 3877 -6563 3923
rect -6517 3877 -6480 3923
rect -6600 3803 -6480 3877
rect -6600 3757 -6563 3803
rect -6517 3757 -6480 3803
rect -6600 3720 -6480 3757
rect -6360 3923 -6240 4020
rect -6360 3877 -6323 3923
rect -6277 3877 -6240 3923
rect -6360 3803 -6240 3877
rect -6360 3757 -6323 3803
rect -6277 3757 -6240 3803
rect -6360 3720 -6240 3757
rect -6120 3923 -6000 4020
rect -6120 3877 -6083 3923
rect -6037 3877 -6000 3923
rect -6120 3803 -6000 3877
rect -6120 3757 -6083 3803
rect -6037 3757 -6000 3803
rect -6120 3720 -6000 3757
<< mvpdiff >>
rect -7080 5603 -6960 5640
rect -7080 5557 -7043 5603
rect -6997 5557 -6960 5603
rect -7080 5483 -6960 5557
rect -7080 5437 -7043 5483
rect -6997 5437 -6960 5483
rect -7080 5363 -6960 5437
rect -7080 5317 -7043 5363
rect -6997 5317 -6960 5363
rect -7080 5280 -6960 5317
rect -6840 5603 -6720 5640
rect -6840 5557 -6803 5603
rect -6757 5557 -6720 5603
rect -6840 5483 -6720 5557
rect -6840 5437 -6803 5483
rect -6757 5437 -6720 5483
rect -6840 5363 -6720 5437
rect -6840 5317 -6803 5363
rect -6757 5317 -6720 5363
rect -6840 5280 -6720 5317
rect -6600 5603 -6480 5640
rect -6600 5557 -6563 5603
rect -6517 5557 -6480 5603
rect -6600 5483 -6480 5557
rect -6600 5437 -6563 5483
rect -6517 5437 -6480 5483
rect -6600 5363 -6480 5437
rect -6600 5317 -6563 5363
rect -6517 5317 -6480 5363
rect -6600 5280 -6480 5317
rect -6360 5603 -6240 5640
rect -6360 5557 -6323 5603
rect -6277 5557 -6240 5603
rect -6360 5483 -6240 5557
rect -6360 5437 -6323 5483
rect -6277 5437 -6240 5483
rect -6360 5363 -6240 5437
rect -6360 5317 -6323 5363
rect -6277 5317 -6240 5363
rect -6360 5280 -6240 5317
rect -6120 5603 -6000 5640
rect -6120 5557 -6083 5603
rect -6037 5557 -6000 5603
rect -6120 5483 -6000 5557
rect -6120 5437 -6083 5483
rect -6037 5437 -6000 5483
rect -6120 5363 -6000 5437
rect -6120 5317 -6083 5363
rect -6037 5317 -6000 5363
rect -6120 5280 -6000 5317
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
rect -6563 -803 -6517 -757
rect -6563 -923 -6517 -877
rect -6563 -1043 -6517 -997
rect -6323 -803 -6277 -757
rect -6323 -923 -6277 -877
rect -6323 -1043 -6277 -997
rect -6083 -803 -6037 -757
rect -6083 -923 -6037 -877
rect -6083 -1043 -6037 -997
<< pdiffc >>
rect -7043 3877 -6997 3923
rect -7043 3757 -6997 3803
rect -6803 3877 -6757 3923
rect -6803 3757 -6757 3803
rect -6563 3877 -6517 3923
rect -6563 3757 -6517 3803
rect -6323 3877 -6277 3923
rect -6323 3757 -6277 3803
rect -6083 3877 -6037 3923
rect -6083 3757 -6037 3803
<< mvpdiffc >>
rect -7043 5557 -6997 5603
rect -7043 5437 -6997 5483
rect -7043 5317 -6997 5363
rect -6803 5557 -6757 5603
rect -6803 5437 -6757 5483
rect -6803 5317 -6757 5363
rect -6563 5557 -6517 5603
rect -6563 5437 -6517 5483
rect -6563 5317 -6517 5363
rect -6323 5557 -6277 5603
rect -6323 5437 -6277 5483
rect -6323 5317 -6277 5363
rect -6083 5557 -6037 5603
rect -6083 5437 -6037 5483
rect -6083 5317 -6037 5363
<< psubdiff >>
rect -7200 6083 -5880 6120
rect -7200 6037 -7163 6083
rect -7117 6037 -7043 6083
rect -6997 6037 -6923 6083
rect -6877 6037 -6803 6083
rect -6757 6037 -6683 6083
rect -6637 6037 -6563 6083
rect -6517 6037 -6443 6083
rect -6397 6037 -6323 6083
rect -6277 6037 -6203 6083
rect -6157 6037 -6083 6083
rect -6037 6037 -5963 6083
rect -5917 6037 -5880 6083
rect -7200 6000 -5880 6037
rect -7200 4643 -5880 4680
rect -7200 4597 -7163 4643
rect -7117 4597 -7043 4643
rect -6997 4597 -6923 4643
rect -6877 4597 -6803 4643
rect -6757 4597 -6683 4643
rect -6637 4597 -6563 4643
rect -6517 4597 -6443 4643
rect -6397 4597 -6323 4643
rect -6277 4597 -6203 4643
rect -6157 4597 -6083 4643
rect -6037 4597 -5963 4643
rect -5917 4597 -5880 4643
rect -7200 4560 -5880 4597
rect -7200 3083 -5880 3120
rect -7200 3037 -7163 3083
rect -7117 3037 -7043 3083
rect -6997 3037 -6923 3083
rect -6877 3037 -6803 3083
rect -6757 3037 -6683 3083
rect -6637 3037 -6563 3083
rect -6517 3037 -6443 3083
rect -6397 3037 -6323 3083
rect -6277 3037 -6203 3083
rect -6157 3037 -6083 3083
rect -6037 3037 -5963 3083
rect -5917 3037 -5880 3083
rect -7200 3000 -5880 3037
rect -7200 2123 -5880 2160
rect -7200 2077 -7163 2123
rect -7117 2077 -7043 2123
rect -6997 2077 -6923 2123
rect -6877 2077 -6803 2123
rect -6757 2077 -6683 2123
rect -6637 2077 -6563 2123
rect -6517 2077 -6443 2123
rect -6397 2077 -6323 2123
rect -6277 2077 -6203 2123
rect -6157 2077 -6083 2123
rect -6037 2077 -5963 2123
rect -5917 2077 -5880 2123
rect -7200 2040 -5880 2077
rect -7200 1643 -5880 1680
rect -7200 1597 -7163 1643
rect -7117 1597 -7043 1643
rect -6997 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6563 1643
rect -6517 1597 -6443 1643
rect -6397 1597 -6323 1643
rect -6277 1597 -6203 1643
rect -6157 1597 -6083 1643
rect -6037 1597 -5963 1643
rect -5917 1597 -5880 1643
rect -7200 1560 -5880 1597
rect -7200 1163 -5880 1200
rect -7200 1117 -7163 1163
rect -7117 1117 -7043 1163
rect -6997 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6563 1163
rect -6517 1117 -6443 1163
rect -6397 1117 -6323 1163
rect -6277 1117 -6203 1163
rect -6157 1117 -6083 1163
rect -6037 1117 -5963 1163
rect -5917 1117 -5880 1163
rect -7200 1080 -5880 1117
rect -7200 683 -5880 720
rect -7200 637 -7163 683
rect -7117 637 -7043 683
rect -6997 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6563 683
rect -6517 637 -6443 683
rect -6397 637 -6323 683
rect -6277 637 -6203 683
rect -6157 637 -6083 683
rect -6037 637 -5963 683
rect -5917 637 -5880 683
rect -7200 600 -5880 637
rect -7200 -277 -5880 -240
rect -7200 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6083 -277
rect -6037 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -360 -5880 -323
rect -7200 -1237 -5880 -1200
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6083 -1237
rect -6037 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1320 -5880 -1283
<< nsubdiff >>
rect -7080 4403 -6000 4440
rect -7080 4357 -7043 4403
rect -6997 4357 -6923 4403
rect -6877 4357 -6803 4403
rect -6757 4357 -6683 4403
rect -6637 4357 -6563 4403
rect -6517 4357 -6443 4403
rect -6397 4357 -6323 4403
rect -6277 4357 -6203 4403
rect -6157 4357 -6083 4403
rect -6037 4357 -6000 4403
rect -7080 4320 -6000 4357
rect -7080 3323 -6000 3360
rect -7080 3277 -7043 3323
rect -6997 3277 -6923 3323
rect -6877 3277 -6803 3323
rect -6757 3277 -6683 3323
rect -6637 3277 -6563 3323
rect -6517 3277 -6443 3323
rect -6397 3277 -6323 3323
rect -6277 3277 -6203 3323
rect -6157 3277 -6083 3323
rect -6037 3277 -6000 3323
rect -7080 3240 -6000 3277
<< mvnsubdiff >>
rect -7080 5843 -6000 5880
rect -7080 5797 -7043 5843
rect -6997 5797 -6923 5843
rect -6877 5797 -6803 5843
rect -6757 5797 -6683 5843
rect -6637 5797 -6563 5843
rect -6517 5797 -6443 5843
rect -6397 5797 -6323 5843
rect -6277 5797 -6203 5843
rect -6157 5797 -6083 5843
rect -6037 5797 -6000 5843
rect -7080 5760 -6000 5797
rect -7080 4883 -6000 4920
rect -7080 4837 -7043 4883
rect -6997 4837 -6923 4883
rect -6877 4837 -6803 4883
rect -6757 4837 -6683 4883
rect -6637 4837 -6563 4883
rect -6517 4837 -6443 4883
rect -6397 4837 -6323 4883
rect -6277 4837 -6203 4883
rect -6157 4837 -6083 4883
rect -6037 4837 -6000 4883
rect -7080 4800 -6000 4837
<< psubdiffcont >>
rect -7163 6037 -7117 6083
rect -7043 6037 -6997 6083
rect -6923 6037 -6877 6083
rect -6803 6037 -6757 6083
rect -6683 6037 -6637 6083
rect -6563 6037 -6517 6083
rect -6443 6037 -6397 6083
rect -6323 6037 -6277 6083
rect -6203 6037 -6157 6083
rect -6083 6037 -6037 6083
rect -5963 6037 -5917 6083
rect -7163 4597 -7117 4643
rect -7043 4597 -6997 4643
rect -6923 4597 -6877 4643
rect -6803 4597 -6757 4643
rect -6683 4597 -6637 4643
rect -6563 4597 -6517 4643
rect -6443 4597 -6397 4643
rect -6323 4597 -6277 4643
rect -6203 4597 -6157 4643
rect -6083 4597 -6037 4643
rect -5963 4597 -5917 4643
rect -7163 3037 -7117 3083
rect -7043 3037 -6997 3083
rect -6923 3037 -6877 3083
rect -6803 3037 -6757 3083
rect -6683 3037 -6637 3083
rect -6563 3037 -6517 3083
rect -6443 3037 -6397 3083
rect -6323 3037 -6277 3083
rect -6203 3037 -6157 3083
rect -6083 3037 -6037 3083
rect -5963 3037 -5917 3083
rect -7163 2077 -7117 2123
rect -7043 2077 -6997 2123
rect -6923 2077 -6877 2123
rect -6803 2077 -6757 2123
rect -6683 2077 -6637 2123
rect -6563 2077 -6517 2123
rect -6443 2077 -6397 2123
rect -6323 2077 -6277 2123
rect -6203 2077 -6157 2123
rect -6083 2077 -6037 2123
rect -5963 2077 -5917 2123
rect -7163 1597 -7117 1643
rect -7043 1597 -6997 1643
rect -6923 1597 -6877 1643
rect -6803 1597 -6757 1643
rect -6683 1597 -6637 1643
rect -6563 1597 -6517 1643
rect -6443 1597 -6397 1643
rect -6323 1597 -6277 1643
rect -6203 1597 -6157 1643
rect -6083 1597 -6037 1643
rect -5963 1597 -5917 1643
rect -7163 1117 -7117 1163
rect -7043 1117 -6997 1163
rect -6923 1117 -6877 1163
rect -6803 1117 -6757 1163
rect -6683 1117 -6637 1163
rect -6563 1117 -6517 1163
rect -6443 1117 -6397 1163
rect -6323 1117 -6277 1163
rect -6203 1117 -6157 1163
rect -6083 1117 -6037 1163
rect -5963 1117 -5917 1163
rect -7163 637 -7117 683
rect -7043 637 -6997 683
rect -6923 637 -6877 683
rect -6803 637 -6757 683
rect -6683 637 -6637 683
rect -6563 637 -6517 683
rect -6443 637 -6397 683
rect -6323 637 -6277 683
rect -6203 637 -6157 683
rect -6083 637 -6037 683
rect -5963 637 -5917 683
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -6563 -323 -6517 -277
rect -6443 -323 -6397 -277
rect -6323 -323 -6277 -277
rect -6203 -323 -6157 -277
rect -6083 -323 -6037 -277
rect -5963 -323 -5917 -277
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
rect -6563 -1283 -6517 -1237
rect -6443 -1283 -6397 -1237
rect -6323 -1283 -6277 -1237
rect -6203 -1283 -6157 -1237
rect -6083 -1283 -6037 -1237
rect -5963 -1283 -5917 -1237
<< nsubdiffcont >>
rect -7043 4357 -6997 4403
rect -6923 4357 -6877 4403
rect -6803 4357 -6757 4403
rect -6683 4357 -6637 4403
rect -6563 4357 -6517 4403
rect -6443 4357 -6397 4403
rect -6323 4357 -6277 4403
rect -6203 4357 -6157 4403
rect -6083 4357 -6037 4403
rect -7043 3277 -6997 3323
rect -6923 3277 -6877 3323
rect -6803 3277 -6757 3323
rect -6683 3277 -6637 3323
rect -6563 3277 -6517 3323
rect -6443 3277 -6397 3323
rect -6323 3277 -6277 3323
rect -6203 3277 -6157 3323
rect -6083 3277 -6037 3323
<< mvnsubdiffcont >>
rect -7043 5797 -6997 5843
rect -6923 5797 -6877 5843
rect -6803 5797 -6757 5843
rect -6683 5797 -6637 5843
rect -6563 5797 -6517 5843
rect -6443 5797 -6397 5843
rect -6323 5797 -6277 5843
rect -6203 5797 -6157 5843
rect -6083 5797 -6037 5843
rect -7043 4837 -6997 4883
rect -6923 4837 -6877 4883
rect -6803 4837 -6757 4883
rect -6683 4837 -6637 4883
rect -6563 4837 -6517 4883
rect -6443 4837 -6397 4883
rect -6323 4837 -6277 4883
rect -6203 4837 -6157 4883
rect -6083 4837 -6037 4883
<< polysilicon >>
rect -6960 5640 -6840 5700
rect -6720 5640 -6600 5700
rect -6480 5640 -6360 5700
rect -6240 5640 -6120 5700
rect -6960 5160 -6840 5280
rect -6720 5160 -6600 5280
rect -6480 5160 -6360 5280
rect -6240 5160 -6120 5280
rect -6960 5123 -6120 5160
rect -6960 5077 -6923 5123
rect -6877 5077 -6803 5123
rect -6757 5077 -6683 5123
rect -6637 5077 -6563 5123
rect -6517 5077 -6443 5123
rect -6397 5077 -6323 5123
rect -6277 5077 -6203 5123
rect -6157 5077 -6120 5123
rect -6960 5040 -6120 5077
rect -6960 4020 -6840 4080
rect -6720 4020 -6600 4080
rect -6480 4020 -6360 4080
rect -6240 4020 -6120 4080
rect -6960 3600 -6840 3720
rect -6720 3600 -6600 3720
rect -6960 3563 -6600 3600
rect -6960 3517 -6923 3563
rect -6877 3517 -6803 3563
rect -6757 3517 -6683 3563
rect -6637 3517 -6600 3563
rect -6960 3480 -6600 3517
rect -6480 3600 -6360 3720
rect -6240 3600 -6120 3720
rect -6480 3563 -6120 3600
rect -6480 3517 -6443 3563
rect -6397 3517 -6323 3563
rect -6277 3517 -6203 3563
rect -6157 3517 -6120 3563
rect -6480 3480 -6120 3517
rect -6960 -517 -6600 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6803 -517
rect -6757 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -600 -6600 -563
rect -6960 -720 -6840 -600
rect -6720 -720 -6600 -600
rect -6480 -517 -6120 -480
rect -6480 -563 -6443 -517
rect -6397 -563 -6323 -517
rect -6277 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -600 -6120 -563
rect -6480 -720 -6360 -600
rect -6240 -720 -6120 -600
rect -6960 -1140 -6840 -1080
rect -6720 -1140 -6600 -1080
rect -6480 -1140 -6360 -1080
rect -6240 -1140 -6120 -1080
<< polycontact >>
rect -6923 5077 -6877 5123
rect -6803 5077 -6757 5123
rect -6683 5077 -6637 5123
rect -6563 5077 -6517 5123
rect -6443 5077 -6397 5123
rect -6323 5077 -6277 5123
rect -6203 5077 -6157 5123
rect -6923 3517 -6877 3563
rect -6803 3517 -6757 3563
rect -6683 3517 -6637 3563
rect -6443 3517 -6397 3563
rect -6323 3517 -6277 3563
rect -6203 3517 -6157 3563
rect -6923 -563 -6877 -517
rect -6803 -563 -6757 -517
rect -6683 -563 -6637 -517
rect -6443 -563 -6397 -517
rect -6323 -563 -6277 -517
rect -6203 -563 -6157 -517
<< metal1 >>
rect -7200 6083 -5880 6120
rect -7200 6037 -7163 6083
rect -7117 6037 -7043 6083
rect -6997 6037 -6923 6083
rect -6877 6037 -6803 6083
rect -6757 6037 -6683 6083
rect -6637 6037 -6563 6083
rect -6517 6037 -6443 6083
rect -6397 6037 -6323 6083
rect -6277 6037 -6203 6083
rect -6157 6037 -6083 6083
rect -6037 6037 -5963 6083
rect -5917 6037 -5880 6083
rect -7200 6000 -5880 6037
rect -7200 5846 -5880 5880
rect -7200 5794 -7046 5846
rect -6994 5843 -6566 5846
rect -6514 5843 -6086 5846
rect -6994 5797 -6923 5843
rect -6877 5797 -6803 5843
rect -6757 5797 -6683 5843
rect -6637 5797 -6566 5843
rect -6514 5797 -6443 5843
rect -6397 5797 -6323 5843
rect -6277 5797 -6203 5843
rect -6157 5797 -6086 5843
rect -6994 5794 -6566 5797
rect -6514 5794 -6086 5797
rect -6034 5794 -5880 5846
rect -7200 5760 -5880 5794
rect -7080 5606 -6960 5640
rect -7080 5554 -7046 5606
rect -6994 5554 -6960 5606
rect -7080 5486 -6960 5554
rect -7080 5434 -7046 5486
rect -6994 5434 -6960 5486
rect -7080 5366 -6960 5434
rect -7080 5314 -7046 5366
rect -6994 5314 -6960 5366
rect -7080 5280 -6960 5314
rect -6840 5606 -6720 5640
rect -6840 5554 -6806 5606
rect -6754 5554 -6720 5606
rect -6840 5486 -6720 5554
rect -6840 5434 -6806 5486
rect -6754 5434 -6720 5486
rect -6840 5366 -6720 5434
rect -6840 5314 -6806 5366
rect -6754 5314 -6720 5366
rect -6840 5280 -6720 5314
rect -6600 5606 -6480 5640
rect -6600 5554 -6566 5606
rect -6514 5554 -6480 5606
rect -6600 5486 -6480 5554
rect -6600 5434 -6566 5486
rect -6514 5434 -6480 5486
rect -6600 5366 -6480 5434
rect -6600 5314 -6566 5366
rect -6514 5314 -6480 5366
rect -6600 5280 -6480 5314
rect -6360 5606 -6240 5640
rect -6360 5554 -6326 5606
rect -6274 5554 -6240 5606
rect -6360 5486 -6240 5554
rect -6360 5434 -6326 5486
rect -6274 5434 -6240 5486
rect -6360 5366 -6240 5434
rect -6360 5314 -6326 5366
rect -6274 5314 -6240 5366
rect -6360 5280 -6240 5314
rect -6120 5606 -6000 5640
rect -6120 5554 -6086 5606
rect -6034 5554 -6000 5606
rect -6120 5486 -6000 5554
rect -6120 5434 -6086 5486
rect -6034 5434 -6000 5486
rect -6120 5366 -6000 5434
rect -6120 5314 -6086 5366
rect -6034 5314 -6000 5366
rect -6120 5280 -6000 5314
rect -6960 5126 -6120 5160
rect -6960 5123 -6566 5126
rect -6514 5123 -6120 5126
rect -6960 5077 -6923 5123
rect -6877 5077 -6803 5123
rect -6757 5077 -6683 5123
rect -6637 5077 -6566 5123
rect -6514 5077 -6443 5123
rect -6397 5077 -6323 5123
rect -6277 5077 -6203 5123
rect -6157 5077 -6120 5123
rect -6960 5074 -6566 5077
rect -6514 5074 -6120 5077
rect -6960 5040 -6120 5074
rect -7200 4883 -5880 4920
rect -7200 4837 -7043 4883
rect -6997 4837 -6923 4883
rect -6877 4837 -6803 4883
rect -6757 4837 -6683 4883
rect -6637 4837 -6563 4883
rect -6517 4837 -6443 4883
rect -6397 4837 -6323 4883
rect -6277 4837 -6203 4883
rect -6157 4837 -6083 4883
rect -6037 4837 -5880 4883
rect -7200 4800 -5880 4837
rect -7200 4643 -5880 4680
rect -7200 4597 -7163 4643
rect -7117 4597 -7043 4643
rect -6997 4597 -6923 4643
rect -6877 4597 -6803 4643
rect -6757 4597 -6683 4643
rect -6637 4597 -6563 4643
rect -6517 4597 -6443 4643
rect -6397 4597 -6323 4643
rect -6277 4597 -6203 4643
rect -6157 4597 -6083 4643
rect -6037 4597 -5963 4643
rect -5917 4597 -5880 4643
rect -7200 4560 -5880 4597
rect -7200 4403 -5880 4440
rect -7200 4357 -7043 4403
rect -6997 4357 -6923 4403
rect -6877 4357 -6803 4403
rect -6757 4357 -6683 4403
rect -6637 4357 -6563 4403
rect -6517 4357 -6443 4403
rect -6397 4357 -6323 4403
rect -6277 4357 -6203 4403
rect -6157 4357 -6083 4403
rect -6037 4357 -5880 4403
rect -7200 4320 -5880 4357
rect -7080 4166 -6000 4200
rect -7080 4114 -7046 4166
rect -6994 4114 -6566 4166
rect -6514 4114 -6086 4166
rect -6034 4114 -6000 4166
rect -7080 4080 -6000 4114
rect -7080 4046 -6960 4080
rect -7080 3994 -7046 4046
rect -6994 3994 -6960 4046
rect -6600 4046 -6480 4080
rect -7080 3926 -6960 3994
rect -7080 3874 -7046 3926
rect -6994 3874 -6960 3926
rect -7080 3806 -6960 3874
rect -7080 3754 -7046 3806
rect -6994 3754 -6960 3806
rect -7080 3720 -6960 3754
rect -6840 3926 -6720 4020
rect -6840 3874 -6806 3926
rect -6754 3874 -6720 3926
rect -6840 3806 -6720 3874
rect -6840 3754 -6806 3806
rect -6754 3754 -6720 3806
rect -6840 3720 -6720 3754
rect -6600 3994 -6566 4046
rect -6514 3994 -6480 4046
rect -6120 4046 -6000 4080
rect -6600 3923 -6480 3994
rect -6600 3877 -6563 3923
rect -6517 3877 -6480 3923
rect -6600 3803 -6480 3877
rect -6600 3757 -6563 3803
rect -6517 3757 -6480 3803
rect -6600 3720 -6480 3757
rect -6360 3926 -6240 4020
rect -6360 3874 -6326 3926
rect -6274 3874 -6240 3926
rect -6360 3806 -6240 3874
rect -6360 3754 -6326 3806
rect -6274 3754 -6240 3806
rect -6360 3720 -6240 3754
rect -6120 3994 -6086 4046
rect -6034 3994 -6000 4046
rect -6120 3926 -6000 3994
rect -6120 3874 -6086 3926
rect -6034 3874 -6000 3926
rect -6120 3806 -6000 3874
rect -6120 3754 -6086 3806
rect -6034 3754 -6000 3806
rect -6120 3720 -6000 3754
rect -6960 3566 -6600 3600
rect -6960 3563 -6806 3566
rect -6754 3563 -6600 3566
rect -6960 3517 -6923 3563
rect -6877 3517 -6806 3563
rect -6754 3517 -6683 3563
rect -6637 3517 -6600 3563
rect -6960 3514 -6806 3517
rect -6754 3514 -6600 3517
rect -6960 3480 -6600 3514
rect -6480 3566 -6120 3600
rect -6480 3563 -6326 3566
rect -6274 3563 -6120 3566
rect -6480 3517 -6443 3563
rect -6397 3517 -6326 3563
rect -6274 3517 -6203 3563
rect -6157 3517 -6120 3563
rect -6480 3514 -6326 3517
rect -6274 3514 -6120 3517
rect -6480 3480 -6120 3514
rect -7200 3326 -5880 3360
rect -7200 3274 -7046 3326
rect -6994 3323 -6086 3326
rect -6994 3277 -6923 3323
rect -6877 3277 -6803 3323
rect -6757 3277 -6683 3323
rect -6637 3277 -6563 3323
rect -6517 3277 -6443 3323
rect -6397 3277 -6323 3323
rect -6277 3277 -6203 3323
rect -6157 3277 -6086 3323
rect -6994 3274 -6086 3277
rect -6034 3274 -5880 3326
rect -7200 3240 -5880 3274
rect -7200 3086 -5880 3120
rect -7200 3083 -7046 3086
rect -6994 3083 -6086 3086
rect -6034 3083 -5880 3086
rect -7200 3037 -7163 3083
rect -7117 3037 -7046 3083
rect -6994 3037 -6923 3083
rect -6877 3037 -6803 3083
rect -6757 3037 -6683 3083
rect -6637 3037 -6563 3083
rect -6517 3037 -6443 3083
rect -6397 3037 -6323 3083
rect -6277 3037 -6203 3083
rect -6157 3037 -6086 3083
rect -6034 3037 -5963 3083
rect -5917 3037 -5880 3083
rect -7200 3034 -7046 3037
rect -6994 3034 -6086 3037
rect -6034 3034 -5880 3037
rect -7200 3000 -5880 3034
rect -7200 2126 -5880 2160
rect -7200 2123 -7046 2126
rect -6994 2123 -6086 2126
rect -6034 2123 -5880 2126
rect -7200 2077 -7163 2123
rect -7117 2077 -7046 2123
rect -6994 2077 -6923 2123
rect -6877 2077 -6803 2123
rect -6757 2077 -6683 2123
rect -6637 2077 -6563 2123
rect -6517 2077 -6443 2123
rect -6397 2077 -6323 2123
rect -6277 2077 -6203 2123
rect -6157 2077 -6086 2123
rect -6034 2077 -5963 2123
rect -5917 2077 -5880 2123
rect -7200 2074 -7046 2077
rect -6994 2074 -6086 2077
rect -6034 2074 -5880 2077
rect -7200 2040 -5880 2074
rect -7200 1646 -5880 1680
rect -7200 1643 -7046 1646
rect -6994 1643 -6086 1646
rect -6034 1643 -5880 1646
rect -7200 1597 -7163 1643
rect -7117 1597 -7046 1643
rect -6994 1597 -6923 1643
rect -6877 1597 -6803 1643
rect -6757 1597 -6683 1643
rect -6637 1597 -6563 1643
rect -6517 1597 -6443 1643
rect -6397 1597 -6323 1643
rect -6277 1597 -6203 1643
rect -6157 1597 -6086 1643
rect -6034 1597 -5963 1643
rect -5917 1597 -5880 1643
rect -7200 1594 -7046 1597
rect -6994 1594 -6086 1597
rect -6034 1594 -5880 1597
rect -7200 1560 -5880 1594
rect -7200 1166 -5880 1200
rect -7200 1163 -7046 1166
rect -6994 1163 -6086 1166
rect -6034 1163 -5880 1166
rect -7200 1117 -7163 1163
rect -7117 1117 -7046 1163
rect -6994 1117 -6923 1163
rect -6877 1117 -6803 1163
rect -6757 1117 -6683 1163
rect -6637 1117 -6563 1163
rect -6517 1117 -6443 1163
rect -6397 1117 -6323 1163
rect -6277 1117 -6203 1163
rect -6157 1117 -6086 1163
rect -6034 1117 -5963 1163
rect -5917 1117 -5880 1163
rect -7200 1114 -7046 1117
rect -6994 1114 -6086 1117
rect -6034 1114 -5880 1117
rect -7200 1080 -5880 1114
rect -7200 686 -5880 720
rect -7200 683 -7046 686
rect -6994 683 -6086 686
rect -6034 683 -5880 686
rect -7200 637 -7163 683
rect -7117 637 -7046 683
rect -6994 637 -6923 683
rect -6877 637 -6803 683
rect -6757 637 -6683 683
rect -6637 637 -6563 683
rect -6517 637 -6443 683
rect -6397 637 -6323 683
rect -6277 637 -6203 683
rect -6157 637 -6086 683
rect -6034 637 -5963 683
rect -5917 637 -5880 683
rect -7200 634 -7046 637
rect -6994 634 -6086 637
rect -6034 634 -5880 637
rect -7200 600 -5880 634
rect -7200 -274 -5880 -240
rect -7200 -277 -7046 -274
rect -6994 -277 -6086 -274
rect -6034 -277 -5880 -274
rect -7200 -323 -7163 -277
rect -7117 -323 -7046 -277
rect -6994 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6086 -277
rect -6034 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -326 -7046 -323
rect -6994 -326 -6086 -323
rect -6034 -326 -5880 -323
rect -7200 -360 -5880 -326
rect -6960 -514 -6600 -480
rect -6960 -517 -6806 -514
rect -6754 -517 -6600 -514
rect -6960 -563 -6923 -517
rect -6877 -563 -6806 -517
rect -6754 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -566 -6806 -563
rect -6754 -566 -6600 -563
rect -6960 -600 -6600 -566
rect -6480 -514 -6120 -480
rect -6480 -517 -6326 -514
rect -6274 -517 -6120 -514
rect -6480 -563 -6443 -517
rect -6397 -563 -6326 -517
rect -6274 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -566 -6326 -563
rect -6274 -566 -6120 -563
rect -6480 -600 -6120 -566
rect -7080 -754 -6960 -720
rect -7080 -806 -7046 -754
rect -6994 -806 -6960 -754
rect -7080 -874 -6960 -806
rect -7080 -926 -7046 -874
rect -6994 -926 -6960 -874
rect -7080 -994 -6960 -926
rect -7080 -1046 -7046 -994
rect -6994 -1046 -6960 -994
rect -7080 -1080 -6960 -1046
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -754 -6480 -720
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -754 -6000 -720
rect -6120 -806 -6086 -754
rect -6034 -806 -6000 -754
rect -6120 -874 -6000 -806
rect -6120 -926 -6086 -874
rect -6034 -926 -6000 -874
rect -6120 -994 -6000 -926
rect -6120 -1046 -6086 -994
rect -6034 -1046 -6000 -994
rect -6120 -1080 -6000 -1046
rect -7200 -1234 -5880 -1200
rect -7200 -1237 -7046 -1234
rect -6994 -1237 -6086 -1234
rect -6034 -1237 -5880 -1234
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7046 -1237
rect -6994 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6086 -1237
rect -6034 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1286 -7046 -1283
rect -6994 -1286 -6086 -1283
rect -6034 -1286 -5880 -1283
rect -7200 -1320 -5880 -1286
<< via1 >>
rect -7046 5843 -6994 5846
rect -6566 5843 -6514 5846
rect -6086 5843 -6034 5846
rect -7046 5797 -7043 5843
rect -7043 5797 -6997 5843
rect -6997 5797 -6994 5843
rect -6566 5797 -6563 5843
rect -6563 5797 -6517 5843
rect -6517 5797 -6514 5843
rect -6086 5797 -6083 5843
rect -6083 5797 -6037 5843
rect -6037 5797 -6034 5843
rect -7046 5794 -6994 5797
rect -6566 5794 -6514 5797
rect -6086 5794 -6034 5797
rect -7046 5603 -6994 5606
rect -7046 5557 -7043 5603
rect -7043 5557 -6997 5603
rect -6997 5557 -6994 5603
rect -7046 5554 -6994 5557
rect -7046 5483 -6994 5486
rect -7046 5437 -7043 5483
rect -7043 5437 -6997 5483
rect -6997 5437 -6994 5483
rect -7046 5434 -6994 5437
rect -7046 5363 -6994 5366
rect -7046 5317 -7043 5363
rect -7043 5317 -6997 5363
rect -6997 5317 -6994 5363
rect -7046 5314 -6994 5317
rect -6806 5603 -6754 5606
rect -6806 5557 -6803 5603
rect -6803 5557 -6757 5603
rect -6757 5557 -6754 5603
rect -6806 5554 -6754 5557
rect -6806 5483 -6754 5486
rect -6806 5437 -6803 5483
rect -6803 5437 -6757 5483
rect -6757 5437 -6754 5483
rect -6806 5434 -6754 5437
rect -6806 5363 -6754 5366
rect -6806 5317 -6803 5363
rect -6803 5317 -6757 5363
rect -6757 5317 -6754 5363
rect -6806 5314 -6754 5317
rect -6566 5603 -6514 5606
rect -6566 5557 -6563 5603
rect -6563 5557 -6517 5603
rect -6517 5557 -6514 5603
rect -6566 5554 -6514 5557
rect -6566 5483 -6514 5486
rect -6566 5437 -6563 5483
rect -6563 5437 -6517 5483
rect -6517 5437 -6514 5483
rect -6566 5434 -6514 5437
rect -6566 5363 -6514 5366
rect -6566 5317 -6563 5363
rect -6563 5317 -6517 5363
rect -6517 5317 -6514 5363
rect -6566 5314 -6514 5317
rect -6326 5603 -6274 5606
rect -6326 5557 -6323 5603
rect -6323 5557 -6277 5603
rect -6277 5557 -6274 5603
rect -6326 5554 -6274 5557
rect -6326 5483 -6274 5486
rect -6326 5437 -6323 5483
rect -6323 5437 -6277 5483
rect -6277 5437 -6274 5483
rect -6326 5434 -6274 5437
rect -6326 5363 -6274 5366
rect -6326 5317 -6323 5363
rect -6323 5317 -6277 5363
rect -6277 5317 -6274 5363
rect -6326 5314 -6274 5317
rect -6086 5603 -6034 5606
rect -6086 5557 -6083 5603
rect -6083 5557 -6037 5603
rect -6037 5557 -6034 5603
rect -6086 5554 -6034 5557
rect -6086 5483 -6034 5486
rect -6086 5437 -6083 5483
rect -6083 5437 -6037 5483
rect -6037 5437 -6034 5483
rect -6086 5434 -6034 5437
rect -6086 5363 -6034 5366
rect -6086 5317 -6083 5363
rect -6083 5317 -6037 5363
rect -6037 5317 -6034 5363
rect -6086 5314 -6034 5317
rect -6566 5123 -6514 5126
rect -6566 5077 -6563 5123
rect -6563 5077 -6517 5123
rect -6517 5077 -6514 5123
rect -6566 5074 -6514 5077
rect -7046 4114 -6994 4166
rect -6566 4114 -6514 4166
rect -6086 4114 -6034 4166
rect -7046 3994 -6994 4046
rect -7046 3923 -6994 3926
rect -7046 3877 -7043 3923
rect -7043 3877 -6997 3923
rect -6997 3877 -6994 3923
rect -7046 3874 -6994 3877
rect -7046 3803 -6994 3806
rect -7046 3757 -7043 3803
rect -7043 3757 -6997 3803
rect -6997 3757 -6994 3803
rect -7046 3754 -6994 3757
rect -6806 3923 -6754 3926
rect -6806 3877 -6803 3923
rect -6803 3877 -6757 3923
rect -6757 3877 -6754 3923
rect -6806 3874 -6754 3877
rect -6806 3803 -6754 3806
rect -6806 3757 -6803 3803
rect -6803 3757 -6757 3803
rect -6757 3757 -6754 3803
rect -6806 3754 -6754 3757
rect -6566 3994 -6514 4046
rect -6326 3923 -6274 3926
rect -6326 3877 -6323 3923
rect -6323 3877 -6277 3923
rect -6277 3877 -6274 3923
rect -6326 3874 -6274 3877
rect -6326 3803 -6274 3806
rect -6326 3757 -6323 3803
rect -6323 3757 -6277 3803
rect -6277 3757 -6274 3803
rect -6326 3754 -6274 3757
rect -6086 3994 -6034 4046
rect -6086 3923 -6034 3926
rect -6086 3877 -6083 3923
rect -6083 3877 -6037 3923
rect -6037 3877 -6034 3923
rect -6086 3874 -6034 3877
rect -6086 3803 -6034 3806
rect -6086 3757 -6083 3803
rect -6083 3757 -6037 3803
rect -6037 3757 -6034 3803
rect -6086 3754 -6034 3757
rect -6806 3563 -6754 3566
rect -6806 3517 -6803 3563
rect -6803 3517 -6757 3563
rect -6757 3517 -6754 3563
rect -6806 3514 -6754 3517
rect -6326 3563 -6274 3566
rect -6326 3517 -6323 3563
rect -6323 3517 -6277 3563
rect -6277 3517 -6274 3563
rect -6326 3514 -6274 3517
rect -7046 3323 -6994 3326
rect -6086 3323 -6034 3326
rect -7046 3277 -7043 3323
rect -7043 3277 -6997 3323
rect -6997 3277 -6994 3323
rect -6086 3277 -6083 3323
rect -6083 3277 -6037 3323
rect -6037 3277 -6034 3323
rect -7046 3274 -6994 3277
rect -6086 3274 -6034 3277
rect -7046 3083 -6994 3086
rect -6086 3083 -6034 3086
rect -7046 3037 -7043 3083
rect -7043 3037 -6997 3083
rect -6997 3037 -6994 3083
rect -6086 3037 -6083 3083
rect -6083 3037 -6037 3083
rect -6037 3037 -6034 3083
rect -7046 3034 -6994 3037
rect -6086 3034 -6034 3037
rect -7046 2123 -6994 2126
rect -6086 2123 -6034 2126
rect -7046 2077 -7043 2123
rect -7043 2077 -6997 2123
rect -6997 2077 -6994 2123
rect -6086 2077 -6083 2123
rect -6083 2077 -6037 2123
rect -6037 2077 -6034 2123
rect -7046 2074 -6994 2077
rect -6086 2074 -6034 2077
rect -7046 1643 -6994 1646
rect -6086 1643 -6034 1646
rect -7046 1597 -7043 1643
rect -7043 1597 -6997 1643
rect -6997 1597 -6994 1643
rect -6086 1597 -6083 1643
rect -6083 1597 -6037 1643
rect -6037 1597 -6034 1643
rect -7046 1594 -6994 1597
rect -6086 1594 -6034 1597
rect -7046 1163 -6994 1166
rect -6086 1163 -6034 1166
rect -7046 1117 -7043 1163
rect -7043 1117 -6997 1163
rect -6997 1117 -6994 1163
rect -6086 1117 -6083 1163
rect -6083 1117 -6037 1163
rect -6037 1117 -6034 1163
rect -7046 1114 -6994 1117
rect -6086 1114 -6034 1117
rect -7046 683 -6994 686
rect -6086 683 -6034 686
rect -7046 637 -7043 683
rect -7043 637 -6997 683
rect -6997 637 -6994 683
rect -6086 637 -6083 683
rect -6083 637 -6037 683
rect -6037 637 -6034 683
rect -7046 634 -6994 637
rect -6086 634 -6034 637
rect -7046 -277 -6994 -274
rect -6086 -277 -6034 -274
rect -7046 -323 -7043 -277
rect -7043 -323 -6997 -277
rect -6997 -323 -6994 -277
rect -6086 -323 -6083 -277
rect -6083 -323 -6037 -277
rect -6037 -323 -6034 -277
rect -7046 -326 -6994 -323
rect -6086 -326 -6034 -323
rect -6806 -517 -6754 -514
rect -6806 -563 -6803 -517
rect -6803 -563 -6757 -517
rect -6757 -563 -6754 -517
rect -6806 -566 -6754 -563
rect -6326 -517 -6274 -514
rect -6326 -563 -6323 -517
rect -6323 -563 -6277 -517
rect -6277 -563 -6274 -517
rect -6326 -566 -6274 -563
rect -7046 -757 -6994 -754
rect -7046 -803 -7043 -757
rect -7043 -803 -6997 -757
rect -6997 -803 -6994 -757
rect -7046 -806 -6994 -803
rect -7046 -877 -6994 -874
rect -7046 -923 -7043 -877
rect -7043 -923 -6997 -877
rect -6997 -923 -6994 -877
rect -7046 -926 -6994 -923
rect -7046 -997 -6994 -994
rect -7046 -1043 -7043 -997
rect -7043 -1043 -6997 -997
rect -6997 -1043 -6994 -997
rect -7046 -1046 -6994 -1043
rect -6566 -757 -6514 -754
rect -6566 -803 -6563 -757
rect -6563 -803 -6517 -757
rect -6517 -803 -6514 -757
rect -6566 -806 -6514 -803
rect -6566 -877 -6514 -874
rect -6566 -923 -6563 -877
rect -6563 -923 -6517 -877
rect -6517 -923 -6514 -877
rect -6566 -926 -6514 -923
rect -6566 -997 -6514 -994
rect -6566 -1043 -6563 -997
rect -6563 -1043 -6517 -997
rect -6517 -1043 -6514 -997
rect -6566 -1046 -6514 -1043
rect -6086 -757 -6034 -754
rect -6086 -803 -6083 -757
rect -6083 -803 -6037 -757
rect -6037 -803 -6034 -757
rect -6086 -806 -6034 -803
rect -6086 -877 -6034 -874
rect -6086 -923 -6083 -877
rect -6083 -923 -6037 -877
rect -6037 -923 -6034 -877
rect -6086 -926 -6034 -923
rect -6086 -997 -6034 -994
rect -6086 -1043 -6083 -997
rect -6083 -1043 -6037 -997
rect -6037 -1043 -6034 -997
rect -6086 -1046 -6034 -1043
rect -7046 -1237 -6994 -1234
rect -6086 -1237 -6034 -1234
rect -7046 -1283 -7043 -1237
rect -7043 -1283 -6997 -1237
rect -6997 -1283 -6994 -1237
rect -6086 -1283 -6083 -1237
rect -6083 -1283 -6037 -1237
rect -6037 -1283 -6034 -1237
rect -7046 -1286 -6994 -1283
rect -6086 -1286 -6034 -1283
<< metal2 >>
rect -7080 5848 -6960 5880
rect -7080 5792 -7048 5848
rect -6992 5792 -6960 5848
rect -7080 5608 -6960 5792
rect -6600 5848 -6480 5880
rect -6600 5792 -6568 5848
rect -6512 5792 -6480 5848
rect -7080 5552 -7048 5608
rect -6992 5552 -6960 5608
rect -7080 5488 -6960 5552
rect -7080 5432 -7048 5488
rect -6992 5432 -6960 5488
rect -7080 5368 -6960 5432
rect -7080 5312 -7048 5368
rect -6992 5312 -6960 5368
rect -7080 5280 -6960 5312
rect -6840 5606 -6720 5640
rect -6840 5554 -6806 5606
rect -6754 5554 -6720 5606
rect -6840 5486 -6720 5554
rect -6840 5434 -6806 5486
rect -6754 5434 -6720 5486
rect -6840 5366 -6720 5434
rect -6840 5314 -6806 5366
rect -6754 5314 -6720 5366
rect -6840 4888 -6720 5314
rect -6600 5608 -6480 5792
rect -6120 5848 -6000 5880
rect -6120 5792 -6088 5848
rect -6032 5792 -6000 5848
rect -6600 5552 -6568 5608
rect -6512 5552 -6480 5608
rect -6600 5488 -6480 5552
rect -6600 5432 -6568 5488
rect -6512 5432 -6480 5488
rect -6600 5368 -6480 5432
rect -6600 5312 -6568 5368
rect -6512 5312 -6480 5368
rect -6600 5280 -6480 5312
rect -6360 5606 -6240 5640
rect -6360 5554 -6326 5606
rect -6274 5554 -6240 5606
rect -6360 5486 -6240 5554
rect -6360 5434 -6326 5486
rect -6274 5434 -6240 5486
rect -6360 5366 -6240 5434
rect -6360 5314 -6326 5366
rect -6274 5314 -6240 5366
rect -6600 5128 -6480 5160
rect -6600 5072 -6568 5128
rect -6512 5072 -6480 5128
rect -6600 5040 -6480 5072
rect -6840 4832 -6808 4888
rect -6752 4832 -6720 4888
rect -7080 4408 -6960 4440
rect -7080 4352 -7048 4408
rect -6992 4352 -6960 4408
rect -7080 4166 -6960 4352
rect -6840 4408 -6720 4832
rect -6360 4888 -6240 5314
rect -6120 5608 -6000 5792
rect -6120 5552 -6088 5608
rect -6032 5552 -6000 5608
rect -6120 5488 -6000 5552
rect -6120 5432 -6088 5488
rect -6032 5432 -6000 5488
rect -6120 5368 -6000 5432
rect -6120 5312 -6088 5368
rect -6032 5312 -6000 5368
rect -6120 5280 -6000 5312
rect -6360 4832 -6328 4888
rect -6272 4832 -6240 4888
rect -6840 4352 -6808 4408
rect -6752 4352 -6720 4408
rect -6840 4320 -6720 4352
rect -6600 4408 -6480 4440
rect -6600 4352 -6568 4408
rect -6512 4352 -6480 4408
rect -7080 4114 -7046 4166
rect -6994 4114 -6960 4166
rect -7080 4046 -6960 4114
rect -7080 3994 -7046 4046
rect -6994 3994 -6960 4046
rect -6600 4166 -6480 4352
rect -6360 4408 -6240 4832
rect -6360 4352 -6328 4408
rect -6272 4352 -6240 4408
rect -6360 4320 -6240 4352
rect -6120 4408 -6000 4440
rect -6120 4352 -6088 4408
rect -6032 4352 -6000 4408
rect -6600 4114 -6566 4166
rect -6514 4114 -6480 4166
rect -6600 4046 -6480 4114
rect -7080 3926 -6960 3994
rect -7080 3874 -7046 3926
rect -6994 3874 -6960 3926
rect -7080 3806 -6960 3874
rect -7080 3754 -7046 3806
rect -6994 3754 -6960 3806
rect -7080 3720 -6960 3754
rect -6840 3926 -6720 4020
rect -6600 3994 -6566 4046
rect -6514 3994 -6480 4046
rect -6120 4166 -6000 4352
rect -6120 4114 -6086 4166
rect -6034 4114 -6000 4166
rect -6120 4046 -6000 4114
rect -6600 3960 -6480 3994
rect -6840 3874 -6806 3926
rect -6754 3874 -6720 3926
rect -6840 3840 -6720 3874
rect -6360 3926 -6240 4020
rect -6360 3874 -6326 3926
rect -6274 3874 -6240 3926
rect -6360 3840 -6240 3874
rect -6840 3806 -6240 3840
rect -6840 3754 -6806 3806
rect -6754 3754 -6326 3806
rect -6274 3754 -6240 3806
rect -6840 3720 -6240 3754
rect -6120 3994 -6086 4046
rect -6034 3994 -6000 4046
rect -6120 3926 -6000 3994
rect -6120 3874 -6086 3926
rect -6034 3874 -6000 3926
rect -6120 3806 -6000 3874
rect -6120 3754 -6086 3806
rect -6034 3754 -6000 3806
rect -6120 3720 -6000 3754
rect -6840 3568 -6720 3600
rect -6840 3512 -6808 3568
rect -6752 3512 -6720 3568
rect -6840 3480 -6720 3512
rect -7080 3328 -6960 3360
rect -7080 3272 -7048 3328
rect -6992 3272 -6960 3328
rect -7080 3240 -6960 3272
rect -7080 3088 -6960 3120
rect -7080 3032 -7048 3088
rect -6992 3032 -6960 3088
rect -7080 2128 -6960 3032
rect -7080 2072 -7048 2128
rect -6992 2072 -6960 2128
rect -7080 1648 -6960 2072
rect -7080 1592 -7048 1648
rect -6992 1592 -6960 1648
rect -7080 1168 -6960 1592
rect -7080 1112 -7048 1168
rect -6992 1112 -6960 1168
rect -7080 688 -6960 1112
rect -7080 632 -7048 688
rect -6992 632 -6960 688
rect -7080 -272 -6960 632
rect -7080 -328 -7048 -272
rect -6992 -328 -6960 -272
rect -7080 -752 -6960 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -7080 -808 -7048 -752
rect -6992 -808 -6960 -752
rect -7080 -872 -6960 -808
rect -7080 -928 -7048 -872
rect -6992 -928 -6960 -872
rect -7080 -992 -6960 -928
rect -7080 -1048 -7048 -992
rect -6992 -1048 -6960 -992
rect -7080 -1232 -6960 -1048
rect -6600 -754 -6480 3720
rect -6360 3568 -6240 3600
rect -6360 3512 -6328 3568
rect -6272 3512 -6240 3568
rect -6360 3480 -6240 3512
rect -6120 3328 -6000 3360
rect -6120 3272 -6088 3328
rect -6032 3272 -6000 3328
rect -6120 3240 -6000 3272
rect -6120 3088 -6000 3120
rect -6120 3032 -6088 3088
rect -6032 3032 -6000 3088
rect -6120 2128 -6000 3032
rect -6120 2072 -6088 2128
rect -6032 2072 -6000 2128
rect -6120 1648 -6000 2072
rect -6120 1592 -6088 1648
rect -6032 1592 -6000 1648
rect -6120 1168 -6000 1592
rect -6120 1112 -6088 1168
rect -6032 1112 -6000 1168
rect -6120 688 -6000 1112
rect -6120 632 -6088 688
rect -6032 632 -6000 688
rect -6120 -272 -6000 632
rect -6120 -328 -6088 -272
rect -6032 -328 -6000 -272
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6120 -752 -6000 -328
rect -6120 -808 -6088 -752
rect -6032 -808 -6000 -752
rect -6120 -872 -6000 -808
rect -6120 -928 -6088 -872
rect -6032 -928 -6000 -872
rect -6120 -992 -6000 -928
rect -6120 -1048 -6088 -992
rect -6032 -1048 -6000 -992
rect -7080 -1288 -7048 -1232
rect -6992 -1288 -6960 -1232
rect -7080 -1320 -6960 -1288
rect -6120 -1232 -6000 -1048
rect -6120 -1288 -6088 -1232
rect -6032 -1288 -6000 -1232
rect -6120 -1320 -6000 -1288
<< via2 >>
rect -7048 5846 -6992 5848
rect -7048 5794 -7046 5846
rect -7046 5794 -6994 5846
rect -6994 5794 -6992 5846
rect -7048 5792 -6992 5794
rect -6568 5846 -6512 5848
rect -6568 5794 -6566 5846
rect -6566 5794 -6514 5846
rect -6514 5794 -6512 5846
rect -6568 5792 -6512 5794
rect -7048 5606 -6992 5608
rect -7048 5554 -7046 5606
rect -7046 5554 -6994 5606
rect -6994 5554 -6992 5606
rect -7048 5552 -6992 5554
rect -7048 5486 -6992 5488
rect -7048 5434 -7046 5486
rect -7046 5434 -6994 5486
rect -6994 5434 -6992 5486
rect -7048 5432 -6992 5434
rect -7048 5366 -6992 5368
rect -7048 5314 -7046 5366
rect -7046 5314 -6994 5366
rect -6994 5314 -6992 5366
rect -7048 5312 -6992 5314
rect -6088 5846 -6032 5848
rect -6088 5794 -6086 5846
rect -6086 5794 -6034 5846
rect -6034 5794 -6032 5846
rect -6088 5792 -6032 5794
rect -6568 5606 -6512 5608
rect -6568 5554 -6566 5606
rect -6566 5554 -6514 5606
rect -6514 5554 -6512 5606
rect -6568 5552 -6512 5554
rect -6568 5486 -6512 5488
rect -6568 5434 -6566 5486
rect -6566 5434 -6514 5486
rect -6514 5434 -6512 5486
rect -6568 5432 -6512 5434
rect -6568 5366 -6512 5368
rect -6568 5314 -6566 5366
rect -6566 5314 -6514 5366
rect -6514 5314 -6512 5366
rect -6568 5312 -6512 5314
rect -6568 5126 -6512 5128
rect -6568 5074 -6566 5126
rect -6566 5074 -6514 5126
rect -6514 5074 -6512 5126
rect -6568 5072 -6512 5074
rect -6808 4832 -6752 4888
rect -7048 4352 -6992 4408
rect -6088 5606 -6032 5608
rect -6088 5554 -6086 5606
rect -6086 5554 -6034 5606
rect -6034 5554 -6032 5606
rect -6088 5552 -6032 5554
rect -6088 5486 -6032 5488
rect -6088 5434 -6086 5486
rect -6086 5434 -6034 5486
rect -6034 5434 -6032 5486
rect -6088 5432 -6032 5434
rect -6088 5366 -6032 5368
rect -6088 5314 -6086 5366
rect -6086 5314 -6034 5366
rect -6034 5314 -6032 5366
rect -6088 5312 -6032 5314
rect -6328 4832 -6272 4888
rect -6808 4352 -6752 4408
rect -6568 4352 -6512 4408
rect -6328 4352 -6272 4408
rect -6088 4352 -6032 4408
rect -6808 3566 -6752 3568
rect -6808 3514 -6806 3566
rect -6806 3514 -6754 3566
rect -6754 3514 -6752 3566
rect -6808 3512 -6752 3514
rect -7048 3326 -6992 3328
rect -7048 3274 -7046 3326
rect -7046 3274 -6994 3326
rect -6994 3274 -6992 3326
rect -7048 3272 -6992 3274
rect -7048 3086 -6992 3088
rect -7048 3034 -7046 3086
rect -7046 3034 -6994 3086
rect -6994 3034 -6992 3086
rect -7048 3032 -6992 3034
rect -7048 2126 -6992 2128
rect -7048 2074 -7046 2126
rect -7046 2074 -6994 2126
rect -6994 2074 -6992 2126
rect -7048 2072 -6992 2074
rect -7048 1646 -6992 1648
rect -7048 1594 -7046 1646
rect -7046 1594 -6994 1646
rect -6994 1594 -6992 1646
rect -7048 1592 -6992 1594
rect -7048 1166 -6992 1168
rect -7048 1114 -7046 1166
rect -7046 1114 -6994 1166
rect -6994 1114 -6992 1166
rect -7048 1112 -6992 1114
rect -7048 686 -6992 688
rect -7048 634 -7046 686
rect -7046 634 -6994 686
rect -6994 634 -6992 686
rect -7048 632 -6992 634
rect -7048 -274 -6992 -272
rect -7048 -326 -7046 -274
rect -7046 -326 -6994 -274
rect -6994 -326 -6992 -274
rect -7048 -328 -6992 -326
rect -6808 -514 -6752 -512
rect -6808 -566 -6806 -514
rect -6806 -566 -6754 -514
rect -6754 -566 -6752 -514
rect -6808 -568 -6752 -566
rect -7048 -754 -6992 -752
rect -7048 -806 -7046 -754
rect -7046 -806 -6994 -754
rect -6994 -806 -6992 -754
rect -7048 -808 -6992 -806
rect -7048 -874 -6992 -872
rect -7048 -926 -7046 -874
rect -7046 -926 -6994 -874
rect -6994 -926 -6992 -874
rect -7048 -928 -6992 -926
rect -7048 -994 -6992 -992
rect -7048 -1046 -7046 -994
rect -7046 -1046 -6994 -994
rect -6994 -1046 -6992 -994
rect -7048 -1048 -6992 -1046
rect -6328 3566 -6272 3568
rect -6328 3514 -6326 3566
rect -6326 3514 -6274 3566
rect -6274 3514 -6272 3566
rect -6328 3512 -6272 3514
rect -6088 3326 -6032 3328
rect -6088 3274 -6086 3326
rect -6086 3274 -6034 3326
rect -6034 3274 -6032 3326
rect -6088 3272 -6032 3274
rect -6088 3086 -6032 3088
rect -6088 3034 -6086 3086
rect -6086 3034 -6034 3086
rect -6034 3034 -6032 3086
rect -6088 3032 -6032 3034
rect -6088 2126 -6032 2128
rect -6088 2074 -6086 2126
rect -6086 2074 -6034 2126
rect -6034 2074 -6032 2126
rect -6088 2072 -6032 2074
rect -6088 1646 -6032 1648
rect -6088 1594 -6086 1646
rect -6086 1594 -6034 1646
rect -6034 1594 -6032 1646
rect -6088 1592 -6032 1594
rect -6088 1166 -6032 1168
rect -6088 1114 -6086 1166
rect -6086 1114 -6034 1166
rect -6034 1114 -6032 1166
rect -6088 1112 -6032 1114
rect -6088 686 -6032 688
rect -6088 634 -6086 686
rect -6086 634 -6034 686
rect -6034 634 -6032 686
rect -6088 632 -6032 634
rect -6088 -274 -6032 -272
rect -6088 -326 -6086 -274
rect -6086 -326 -6034 -274
rect -6034 -326 -6032 -274
rect -6088 -328 -6032 -326
rect -6328 -514 -6272 -512
rect -6328 -566 -6326 -514
rect -6326 -566 -6274 -514
rect -6274 -566 -6272 -514
rect -6328 -568 -6272 -566
rect -6088 -754 -6032 -752
rect -6088 -806 -6086 -754
rect -6086 -806 -6034 -754
rect -6034 -806 -6032 -754
rect -6088 -808 -6032 -806
rect -6088 -874 -6032 -872
rect -6088 -926 -6086 -874
rect -6086 -926 -6034 -874
rect -6034 -926 -6032 -874
rect -6088 -928 -6032 -926
rect -6088 -994 -6032 -992
rect -6088 -1046 -6086 -994
rect -6086 -1046 -6034 -994
rect -6034 -1046 -6032 -994
rect -6088 -1048 -6032 -1046
rect -7048 -1234 -6992 -1232
rect -7048 -1286 -7046 -1234
rect -7046 -1286 -6994 -1234
rect -6994 -1286 -6992 -1234
rect -7048 -1288 -6992 -1286
rect -6088 -1234 -6032 -1232
rect -6088 -1286 -6086 -1234
rect -6086 -1286 -6034 -1234
rect -6034 -1286 -6032 -1234
rect -6088 -1288 -6032 -1286
<< metal3 >>
rect -7200 5848 -5880 5880
rect -7200 5792 -7048 5848
rect -6992 5792 -6568 5848
rect -6512 5792 -6088 5848
rect -6032 5792 -5880 5848
rect -7200 5608 -5880 5792
rect -7200 5552 -7048 5608
rect -6992 5552 -6568 5608
rect -6512 5552 -6088 5608
rect -6032 5552 -5880 5608
rect -7200 5488 -5880 5552
rect -7200 5432 -7048 5488
rect -6992 5432 -6568 5488
rect -6512 5432 -6088 5488
rect -6032 5432 -5880 5488
rect -7200 5368 -5880 5432
rect -7200 5312 -7048 5368
rect -6992 5312 -6568 5368
rect -6512 5312 -6088 5368
rect -6032 5312 -5880 5368
rect -7200 5280 -5880 5312
rect -6600 5128 -6480 5160
rect -6600 5072 -6568 5128
rect -6512 5072 -6480 5128
rect -6600 5040 -6480 5072
rect -7200 4888 -5880 4920
rect -7200 4832 -6808 4888
rect -6752 4832 -6328 4888
rect -6272 4832 -5880 4888
rect -7200 4740 -5880 4832
rect -7200 4648 -5880 4680
rect -7200 4592 -6568 4648
rect -6512 4592 -5880 4648
rect -7200 4560 -5880 4592
rect -7200 4408 -5880 4500
rect -7200 4352 -7048 4408
rect -6992 4352 -6808 4408
rect -6752 4352 -6568 4408
rect -6512 4352 -6328 4408
rect -6272 4352 -6088 4408
rect -6032 4352 -5880 4408
rect -7200 4320 -5880 4352
rect -6840 3568 -6720 3600
rect -6840 3512 -6808 3568
rect -6752 3512 -6720 3568
rect -6840 3480 -6720 3512
rect -6360 3568 -6240 3600
rect -6360 3512 -6328 3568
rect -6272 3512 -6240 3568
rect -6360 3480 -6240 3512
rect -7200 3328 -5880 3360
rect -7200 3272 -7048 3328
rect -6992 3272 -6088 3328
rect -6032 3272 -5880 3328
rect -7200 3240 -5880 3272
rect -7200 3088 -5880 3120
rect -7200 3032 -7048 3088
rect -6992 3032 -6088 3088
rect -6032 3032 -5880 3088
rect -7200 3000 -5880 3032
rect -7200 2280 -5880 2880
rect -7200 2128 -5880 2160
rect -7200 2072 -7048 2128
rect -6992 2072 -6088 2128
rect -6032 2072 -5880 2128
rect -7200 2040 -5880 2072
rect -7200 1800 -5880 1920
rect -7200 1648 -5880 1680
rect -7200 1592 -7048 1648
rect -6992 1592 -6088 1648
rect -6032 1592 -5880 1648
rect -7200 1560 -5880 1592
rect -7200 1320 -5880 1440
rect -7200 1168 -5880 1200
rect -7200 1112 -7048 1168
rect -6992 1112 -6088 1168
rect -6032 1112 -5880 1168
rect -7200 1080 -5880 1112
rect -7200 840 -5880 960
rect -7200 688 -5880 720
rect -7200 632 -7048 688
rect -6992 632 -6088 688
rect -6032 632 -5880 688
rect -7200 600 -5880 632
rect -7200 -120 -5880 480
rect -7200 -272 -5880 -240
rect -7200 -328 -7048 -272
rect -6992 -328 -6088 -272
rect -6032 -328 -5880 -272
rect -7200 -360 -5880 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -7200 -752 -5880 -720
rect -7200 -808 -7048 -752
rect -6992 -808 -6088 -752
rect -6032 -808 -5880 -752
rect -7200 -872 -5880 -808
rect -7200 -928 -7048 -872
rect -6992 -928 -6088 -872
rect -6032 -928 -5880 -872
rect -7200 -992 -5880 -928
rect -7200 -1048 -7048 -992
rect -6992 -1048 -6088 -992
rect -6032 -1048 -5880 -992
rect -7200 -1232 -5880 -1048
rect -7200 -1288 -7048 -1232
rect -6992 -1288 -6088 -1232
rect -6032 -1288 -5880 -1232
rect -7200 -1320 -5880 -1288
<< via3 >>
rect -6568 5072 -6512 5128
rect -6808 4832 -6752 4888
rect -6328 4832 -6272 4888
rect -6568 4592 -6512 4648
rect -7048 4352 -6992 4408
rect -6808 4352 -6752 4408
rect -6328 4352 -6272 4408
rect -6088 4352 -6032 4408
rect -6808 3512 -6752 3568
rect -6328 3512 -6272 3568
rect -6808 -568 -6752 -512
rect -6328 -568 -6272 -512
<< metal4 >>
rect -6600 5128 -6480 5160
rect -6600 5072 -6568 5128
rect -6512 5072 -6480 5128
rect -6840 4888 -6720 4920
rect -6840 4832 -6808 4888
rect -6752 4832 -6720 4888
rect -7080 4408 -6960 4440
rect -7080 4352 -7048 4408
rect -6992 4352 -6960 4408
rect -7080 4320 -6960 4352
rect -6840 4408 -6720 4832
rect -6600 4648 -6480 5072
rect -6600 4592 -6568 4648
rect -6512 4592 -6480 4648
rect -6600 4560 -6480 4592
rect -6360 4888 -6240 4920
rect -6360 4832 -6328 4888
rect -6272 4832 -6240 4888
rect -6840 4352 -6808 4408
rect -6752 4352 -6720 4408
rect -6840 4320 -6720 4352
rect -6360 4408 -6240 4832
rect -6360 4352 -6328 4408
rect -6272 4352 -6240 4408
rect -6360 4320 -6240 4352
rect -6120 4408 -6000 4440
rect -6120 4352 -6088 4408
rect -6032 4352 -6000 4408
rect -6120 4320 -6000 4352
rect -6840 3568 -6720 3600
rect -6840 3512 -6808 3568
rect -6752 3512 -6720 3568
rect -6840 3360 -6720 3512
rect -7080 3240 -6720 3360
rect -6840 -512 -6720 3240
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 3568 -6240 3600
rect -6360 3512 -6328 3568
rect -6272 3512 -6240 3568
rect -6360 3360 -6240 3512
rect -6360 3240 -6000 3360
rect -6360 -512 -6240 3240
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
<< labels >>
rlabel metal1 s -6780 -900 -6780 -900 4 d1
rlabel metal1 s -6300 -900 -6300 -900 4 d2
rlabel metal1 s -6540 6060 -6540 6060 4 vss
rlabel metal1 s -6540 4620 -6540 4620 4 vss
rlabel metal4 s -6840 -120 -6720 2400 4 inl
port 1 nsew
rlabel metal4 s -6360 -120 -6240 2400 4 inr
port 2 nsew
rlabel metal2 s -6600 -120 -6480 2400 4 out
port 3 nsew
rlabel metal3 s -7200 5280 -5880 5880 4 vdd
port 4 nsew
rlabel metal3 s -7200 4560 -5880 4680 4 gp
port 5 nsew
rlabel metal3 s -7200 4740 -7080 4920 4 vreg
port 6 nsew
rlabel metal3 s -7200 2280 -5880 2880 4 op
port 7 nsew
rlabel metal3 s -7200 1800 -5880 1920 4 im
port 8 nsew
rlabel metal3 s -7200 840 -5880 960 4 ip
port 9 nsew
rlabel metal3 s -7200 -120 -5880 480 4 om
port 10 nsew
rlabel metal3 s -7200 -1320 -5880 -720 4 gnd
port 11 nsew
<< end >>
