* Amplifier open-loop DC testbench

* Include GF180MCU device models
.include "../../../gf180mcuC/libs.tech/ngspice/design.ngspice"
.lib "../../../gf180mcuC/libs.tech/ngspice/sm141064.ngspice" typical

.include "inv.spice"
.include "../magic/inv.spice"

.param pVDH = 5.0
.param pVDX = 3.3
.param pIB  = 20.0u

VDH vdh 0 dc {pVDH}
VDX vdx 0 dc {pVDX}
VSS vss 0 0
ECM cm vss vdx vss 0.5

vin in cm dc 0 ac 1

*ib vdd ib {pIB}
xb ib      vdh vdh bp  vdx vss inv_bias
x0 in  out vdh vdh bp  vdx vss inv0
evdq vdq vss vdx vss 1
xq q   q   vdh vdh bp  vdq vss inv0
vo out cm
.param dx = 1.5
.dc vin {-dx} {dx} {dx/1001}
.option gmin = 1e-15
.control	
	alter vdx dc=3.0
	dc vin -1.5 1.5 1m
		
	let vi = in-cm
	let io = i(vo)
	let gm = abs(deriv(io))
	
	meas dc iq  find i(evdq) at=0
	meas dc io0 find io at=0
	meas dc gm0 find gm at=0
	let ioN = i(vo)/gm0
	let gmN = gm/gm0

	wrdata ../data/inv_gm_vdd30.txt io gm ioN gmN

	alter vdx dc=2.4
	dc vin -1.2 1.2 1m

	let vi = in-cm
	let io = i(vo)
	let gm = abs(deriv(io))

	meas dc iq  find i(evdq) at=0	
	meas dc io0 find io at=0
	meas dc gm0 find gm at=0
	let ioN = i(vo)/gm0
	let gmN = gm/gm0

	wrdata ../data/inv_gm_vdd24.txt io gm ioN gmN

	alter vdx dc=1.8
	dc vin -0.9 0.9 1m

	let vi = in-cm
	let io = i(vo)
	let gm = abs(deriv(io))

	meas dc iq  find i(evdq) at=0	
	meas dc io0 find io at=0
	meas dc gm0 find gm at=0
	let ioN = i(vo)/gm0
	let gmN = gm/gm0

	wrdata ../data/inv_gm_vdd18.txt io gm ioN gmN

	plot dc1.io dc2.io dc3.io
	plot dc1.gm dc2.gm dc3.gm
	
	plot dc1.ion dc2.ion dc3.ion
	plot dc1.gmn dc2.gmn dc3.gmn



.endc

.end
