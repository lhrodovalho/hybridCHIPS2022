magic
tech gf180mcuC
magscale 1 10
timestamp 1665184495
<< nwell >>
rect -7200 5700 -5880 6900
rect -7200 4140 -5880 5460
<< nmos >>
rect -6960 -1080 -6840 -720
rect -6720 -1080 -6600 -720
rect -6480 -1080 -6360 -720
rect -6240 -1080 -6120 -720
<< pmos >>
rect -6960 4680 -6840 4980
rect -6720 4680 -6600 4980
rect -6480 4680 -6360 4980
rect -6240 4680 -6120 4980
<< mvpmos >>
rect -6960 6240 -6840 6600
rect -6720 6240 -6600 6600
rect -6480 6240 -6360 6600
rect -6240 6240 -6120 6600
<< ndiff >>
rect -7080 -757 -6960 -720
rect -7080 -803 -7043 -757
rect -6997 -803 -6960 -757
rect -7080 -877 -6960 -803
rect -7080 -923 -7043 -877
rect -6997 -923 -6960 -877
rect -7080 -997 -6960 -923
rect -7080 -1043 -7043 -997
rect -6997 -1043 -6960 -997
rect -7080 -1080 -6960 -1043
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -757 -6480 -720
rect -6600 -803 -6563 -757
rect -6517 -803 -6480 -757
rect -6600 -877 -6480 -803
rect -6600 -923 -6563 -877
rect -6517 -923 -6480 -877
rect -6600 -997 -6480 -923
rect -6600 -1043 -6563 -997
rect -6517 -1043 -6480 -997
rect -6600 -1080 -6480 -1043
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -757 -6000 -720
rect -6120 -803 -6083 -757
rect -6037 -803 -6000 -757
rect -6120 -877 -6000 -803
rect -6120 -923 -6083 -877
rect -6037 -923 -6000 -877
rect -6120 -997 -6000 -923
rect -6120 -1043 -6083 -997
rect -6037 -1043 -6000 -997
rect -6120 -1080 -6000 -1043
<< pdiff >>
rect -7080 4883 -6960 4980
rect -7080 4837 -7043 4883
rect -6997 4837 -6960 4883
rect -7080 4763 -6960 4837
rect -7080 4717 -7043 4763
rect -6997 4717 -6960 4763
rect -7080 4680 -6960 4717
rect -6840 4883 -6720 4980
rect -6840 4837 -6803 4883
rect -6757 4837 -6720 4883
rect -6840 4763 -6720 4837
rect -6840 4717 -6803 4763
rect -6757 4717 -6720 4763
rect -6840 4680 -6720 4717
rect -6600 4883 -6480 4980
rect -6600 4837 -6563 4883
rect -6517 4837 -6480 4883
rect -6600 4763 -6480 4837
rect -6600 4717 -6563 4763
rect -6517 4717 -6480 4763
rect -6600 4680 -6480 4717
rect -6360 4883 -6240 4980
rect -6360 4837 -6323 4883
rect -6277 4837 -6240 4883
rect -6360 4763 -6240 4837
rect -6360 4717 -6323 4763
rect -6277 4717 -6240 4763
rect -6360 4680 -6240 4717
rect -6120 4883 -6000 4980
rect -6120 4837 -6083 4883
rect -6037 4837 -6000 4883
rect -6120 4763 -6000 4837
rect -6120 4717 -6083 4763
rect -6037 4717 -6000 4763
rect -6120 4680 -6000 4717
<< mvpdiff >>
rect -7080 6563 -6960 6600
rect -7080 6517 -7043 6563
rect -6997 6517 -6960 6563
rect -7080 6443 -6960 6517
rect -7080 6397 -7043 6443
rect -6997 6397 -6960 6443
rect -7080 6323 -6960 6397
rect -7080 6277 -7043 6323
rect -6997 6277 -6960 6323
rect -7080 6240 -6960 6277
rect -6840 6563 -6720 6600
rect -6840 6517 -6803 6563
rect -6757 6517 -6720 6563
rect -6840 6443 -6720 6517
rect -6840 6397 -6803 6443
rect -6757 6397 -6720 6443
rect -6840 6323 -6720 6397
rect -6840 6277 -6803 6323
rect -6757 6277 -6720 6323
rect -6840 6240 -6720 6277
rect -6600 6563 -6480 6600
rect -6600 6517 -6563 6563
rect -6517 6517 -6480 6563
rect -6600 6443 -6480 6517
rect -6600 6397 -6563 6443
rect -6517 6397 -6480 6443
rect -6600 6323 -6480 6397
rect -6600 6277 -6563 6323
rect -6517 6277 -6480 6323
rect -6600 6240 -6480 6277
rect -6360 6563 -6240 6600
rect -6360 6517 -6323 6563
rect -6277 6517 -6240 6563
rect -6360 6443 -6240 6517
rect -6360 6397 -6323 6443
rect -6277 6397 -6240 6443
rect -6360 6323 -6240 6397
rect -6360 6277 -6323 6323
rect -6277 6277 -6240 6323
rect -6360 6240 -6240 6277
rect -6120 6563 -6000 6600
rect -6120 6517 -6083 6563
rect -6037 6517 -6000 6563
rect -6120 6443 -6000 6517
rect -6120 6397 -6083 6443
rect -6037 6397 -6000 6443
rect -6120 6323 -6000 6397
rect -6120 6277 -6083 6323
rect -6037 6277 -6000 6323
rect -6120 6240 -6000 6277
<< ndiffc >>
rect -7043 -803 -6997 -757
rect -7043 -923 -6997 -877
rect -7043 -1043 -6997 -997
rect -6803 -803 -6757 -757
rect -6803 -923 -6757 -877
rect -6803 -1043 -6757 -997
rect -6563 -803 -6517 -757
rect -6563 -923 -6517 -877
rect -6563 -1043 -6517 -997
rect -6323 -803 -6277 -757
rect -6323 -923 -6277 -877
rect -6323 -1043 -6277 -997
rect -6083 -803 -6037 -757
rect -6083 -923 -6037 -877
rect -6083 -1043 -6037 -997
<< pdiffc >>
rect -7043 4837 -6997 4883
rect -7043 4717 -6997 4763
rect -6803 4837 -6757 4883
rect -6803 4717 -6757 4763
rect -6563 4837 -6517 4883
rect -6563 4717 -6517 4763
rect -6323 4837 -6277 4883
rect -6323 4717 -6277 4763
rect -6083 4837 -6037 4883
rect -6083 4717 -6037 4763
<< mvpdiffc >>
rect -7043 6517 -6997 6563
rect -7043 6397 -6997 6443
rect -7043 6277 -6997 6323
rect -6803 6517 -6757 6563
rect -6803 6397 -6757 6443
rect -6803 6277 -6757 6323
rect -6563 6517 -6517 6563
rect -6563 6397 -6517 6443
rect -6563 6277 -6517 6323
rect -6323 6517 -6277 6563
rect -6323 6397 -6277 6443
rect -6323 6277 -6277 6323
rect -6083 6517 -6037 6563
rect -6083 6397 -6037 6443
rect -6083 6277 -6037 6323
<< psubdiff >>
rect -7200 7043 -5880 7080
rect -7200 6997 -7163 7043
rect -7117 6997 -7043 7043
rect -6997 6997 -6923 7043
rect -6877 6997 -6803 7043
rect -6757 6997 -6683 7043
rect -6637 6997 -6563 7043
rect -6517 6997 -6443 7043
rect -6397 6997 -6323 7043
rect -6277 6997 -6203 7043
rect -6157 6997 -6083 7043
rect -6037 6997 -5963 7043
rect -5917 6997 -5880 7043
rect -7200 6960 -5880 6997
rect -7200 5603 -5880 5640
rect -7200 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6563 5603
rect -6517 5557 -6443 5603
rect -6397 5557 -6323 5603
rect -6277 5557 -6203 5603
rect -6157 5557 -6083 5603
rect -6037 5557 -5963 5603
rect -5917 5557 -5880 5603
rect -7200 5520 -5880 5557
rect -7200 4043 -5880 4080
rect -7200 3997 -7163 4043
rect -7117 3997 -7043 4043
rect -6997 3997 -6923 4043
rect -6877 3997 -6803 4043
rect -6757 3997 -6683 4043
rect -6637 3997 -6563 4043
rect -6517 3997 -6443 4043
rect -6397 3997 -6323 4043
rect -6277 3997 -6203 4043
rect -6157 3997 -6083 4043
rect -6037 3997 -5963 4043
rect -5917 3997 -5880 4043
rect -7200 3960 -5880 3997
rect -7200 2843 -5880 2880
rect -7200 2797 -7163 2843
rect -7117 2797 -7043 2843
rect -6997 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6683 2843
rect -6637 2797 -6563 2843
rect -6517 2797 -6443 2843
rect -6397 2797 -6323 2843
rect -6277 2797 -6203 2843
rect -6157 2797 -6083 2843
rect -6037 2797 -5963 2843
rect -5917 2797 -5880 2843
rect -7200 2760 -5880 2797
rect -7200 2363 -5880 2400
rect -7200 2317 -7163 2363
rect -7117 2317 -7043 2363
rect -6997 2317 -6923 2363
rect -6877 2317 -6803 2363
rect -6757 2317 -6683 2363
rect -6637 2317 -6563 2363
rect -6517 2317 -6443 2363
rect -6397 2317 -6323 2363
rect -6277 2317 -6203 2363
rect -6157 2317 -6083 2363
rect -6037 2317 -5963 2363
rect -5917 2317 -5880 2363
rect -7200 2280 -5880 2317
rect -7200 1883 -5880 1920
rect -7200 1837 -7163 1883
rect -7117 1837 -7043 1883
rect -6997 1837 -6923 1883
rect -6877 1837 -6803 1883
rect -6757 1837 -6683 1883
rect -6637 1837 -6563 1883
rect -6517 1837 -6443 1883
rect -6397 1837 -6323 1883
rect -6277 1837 -6203 1883
rect -6157 1837 -6083 1883
rect -6037 1837 -5963 1883
rect -5917 1837 -5880 1883
rect -7200 1800 -5880 1837
rect -7200 1403 -5880 1440
rect -7200 1357 -7163 1403
rect -7117 1357 -7043 1403
rect -6997 1357 -6923 1403
rect -6877 1357 -6803 1403
rect -6757 1357 -6683 1403
rect -6637 1357 -6563 1403
rect -6517 1357 -6443 1403
rect -6397 1357 -6323 1403
rect -6277 1357 -6203 1403
rect -6157 1357 -6083 1403
rect -6037 1357 -5963 1403
rect -5917 1357 -5880 1403
rect -7200 1320 -5880 1357
rect -7200 923 -5880 960
rect -7200 877 -7163 923
rect -7117 877 -7043 923
rect -6997 877 -6923 923
rect -6877 877 -6803 923
rect -6757 877 -6683 923
rect -6637 877 -6563 923
rect -6517 877 -6443 923
rect -6397 877 -6323 923
rect -6277 877 -6203 923
rect -6157 877 -6083 923
rect -6037 877 -5963 923
rect -5917 877 -5880 923
rect -7200 840 -5880 877
rect -7200 -277 -5880 -240
rect -7200 -323 -7163 -277
rect -7117 -323 -7043 -277
rect -6997 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6083 -277
rect -6037 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -360 -5880 -323
rect -7200 -1237 -5880 -1200
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7043 -1237
rect -6997 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6083 -1237
rect -6037 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1320 -5880 -1283
<< nsubdiff >>
rect -7080 5363 -6000 5400
rect -7080 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6683 5363
rect -6637 5317 -6563 5363
rect -6517 5317 -6443 5363
rect -6397 5317 -6323 5363
rect -6277 5317 -6203 5363
rect -6157 5317 -6083 5363
rect -6037 5317 -6000 5363
rect -7080 5280 -6000 5317
rect -7080 4283 -6000 4320
rect -7080 4237 -7043 4283
rect -6997 4237 -6923 4283
rect -6877 4237 -6803 4283
rect -6757 4237 -6683 4283
rect -6637 4237 -6563 4283
rect -6517 4237 -6443 4283
rect -6397 4237 -6323 4283
rect -6277 4237 -6203 4283
rect -6157 4237 -6083 4283
rect -6037 4237 -6000 4283
rect -7080 4200 -6000 4237
<< mvnsubdiff >>
rect -7080 6803 -6000 6840
rect -7080 6757 -7043 6803
rect -6997 6757 -6923 6803
rect -6877 6757 -6803 6803
rect -6757 6757 -6683 6803
rect -6637 6757 -6563 6803
rect -6517 6757 -6443 6803
rect -6397 6757 -6323 6803
rect -6277 6757 -6203 6803
rect -6157 6757 -6083 6803
rect -6037 6757 -6000 6803
rect -7080 6720 -6000 6757
rect -7080 5843 -6000 5880
rect -7080 5797 -7043 5843
rect -6997 5797 -6923 5843
rect -6877 5797 -6803 5843
rect -6757 5797 -6683 5843
rect -6637 5797 -6563 5843
rect -6517 5797 -6443 5843
rect -6397 5797 -6323 5843
rect -6277 5797 -6203 5843
rect -6157 5797 -6083 5843
rect -6037 5797 -6000 5843
rect -7080 5760 -6000 5797
<< psubdiffcont >>
rect -7163 6997 -7117 7043
rect -7043 6997 -6997 7043
rect -6923 6997 -6877 7043
rect -6803 6997 -6757 7043
rect -6683 6997 -6637 7043
rect -6563 6997 -6517 7043
rect -6443 6997 -6397 7043
rect -6323 6997 -6277 7043
rect -6203 6997 -6157 7043
rect -6083 6997 -6037 7043
rect -5963 6997 -5917 7043
rect -7163 5557 -7117 5603
rect -7043 5557 -6997 5603
rect -6923 5557 -6877 5603
rect -6803 5557 -6757 5603
rect -6683 5557 -6637 5603
rect -6563 5557 -6517 5603
rect -6443 5557 -6397 5603
rect -6323 5557 -6277 5603
rect -6203 5557 -6157 5603
rect -6083 5557 -6037 5603
rect -5963 5557 -5917 5603
rect -7163 3997 -7117 4043
rect -7043 3997 -6997 4043
rect -6923 3997 -6877 4043
rect -6803 3997 -6757 4043
rect -6683 3997 -6637 4043
rect -6563 3997 -6517 4043
rect -6443 3997 -6397 4043
rect -6323 3997 -6277 4043
rect -6203 3997 -6157 4043
rect -6083 3997 -6037 4043
rect -5963 3997 -5917 4043
rect -7163 2797 -7117 2843
rect -7043 2797 -6997 2843
rect -6923 2797 -6877 2843
rect -6803 2797 -6757 2843
rect -6683 2797 -6637 2843
rect -6563 2797 -6517 2843
rect -6443 2797 -6397 2843
rect -6323 2797 -6277 2843
rect -6203 2797 -6157 2843
rect -6083 2797 -6037 2843
rect -5963 2797 -5917 2843
rect -7163 2317 -7117 2363
rect -7043 2317 -6997 2363
rect -6923 2317 -6877 2363
rect -6803 2317 -6757 2363
rect -6683 2317 -6637 2363
rect -6563 2317 -6517 2363
rect -6443 2317 -6397 2363
rect -6323 2317 -6277 2363
rect -6203 2317 -6157 2363
rect -6083 2317 -6037 2363
rect -5963 2317 -5917 2363
rect -7163 1837 -7117 1883
rect -7043 1837 -6997 1883
rect -6923 1837 -6877 1883
rect -6803 1837 -6757 1883
rect -6683 1837 -6637 1883
rect -6563 1837 -6517 1883
rect -6443 1837 -6397 1883
rect -6323 1837 -6277 1883
rect -6203 1837 -6157 1883
rect -6083 1837 -6037 1883
rect -5963 1837 -5917 1883
rect -7163 1357 -7117 1403
rect -7043 1357 -6997 1403
rect -6923 1357 -6877 1403
rect -6803 1357 -6757 1403
rect -6683 1357 -6637 1403
rect -6563 1357 -6517 1403
rect -6443 1357 -6397 1403
rect -6323 1357 -6277 1403
rect -6203 1357 -6157 1403
rect -6083 1357 -6037 1403
rect -5963 1357 -5917 1403
rect -7163 877 -7117 923
rect -7043 877 -6997 923
rect -6923 877 -6877 923
rect -6803 877 -6757 923
rect -6683 877 -6637 923
rect -6563 877 -6517 923
rect -6443 877 -6397 923
rect -6323 877 -6277 923
rect -6203 877 -6157 923
rect -6083 877 -6037 923
rect -5963 877 -5917 923
rect -7163 -323 -7117 -277
rect -7043 -323 -6997 -277
rect -6923 -323 -6877 -277
rect -6803 -323 -6757 -277
rect -6683 -323 -6637 -277
rect -6563 -323 -6517 -277
rect -6443 -323 -6397 -277
rect -6323 -323 -6277 -277
rect -6203 -323 -6157 -277
rect -6083 -323 -6037 -277
rect -5963 -323 -5917 -277
rect -7163 -1283 -7117 -1237
rect -7043 -1283 -6997 -1237
rect -6923 -1283 -6877 -1237
rect -6803 -1283 -6757 -1237
rect -6683 -1283 -6637 -1237
rect -6563 -1283 -6517 -1237
rect -6443 -1283 -6397 -1237
rect -6323 -1283 -6277 -1237
rect -6203 -1283 -6157 -1237
rect -6083 -1283 -6037 -1237
rect -5963 -1283 -5917 -1237
<< nsubdiffcont >>
rect -7043 5317 -6997 5363
rect -6923 5317 -6877 5363
rect -6803 5317 -6757 5363
rect -6683 5317 -6637 5363
rect -6563 5317 -6517 5363
rect -6443 5317 -6397 5363
rect -6323 5317 -6277 5363
rect -6203 5317 -6157 5363
rect -6083 5317 -6037 5363
rect -7043 4237 -6997 4283
rect -6923 4237 -6877 4283
rect -6803 4237 -6757 4283
rect -6683 4237 -6637 4283
rect -6563 4237 -6517 4283
rect -6443 4237 -6397 4283
rect -6323 4237 -6277 4283
rect -6203 4237 -6157 4283
rect -6083 4237 -6037 4283
<< mvnsubdiffcont >>
rect -7043 6757 -6997 6803
rect -6923 6757 -6877 6803
rect -6803 6757 -6757 6803
rect -6683 6757 -6637 6803
rect -6563 6757 -6517 6803
rect -6443 6757 -6397 6803
rect -6323 6757 -6277 6803
rect -6203 6757 -6157 6803
rect -6083 6757 -6037 6803
rect -7043 5797 -6997 5843
rect -6923 5797 -6877 5843
rect -6803 5797 -6757 5843
rect -6683 5797 -6637 5843
rect -6563 5797 -6517 5843
rect -6443 5797 -6397 5843
rect -6323 5797 -6277 5843
rect -6203 5797 -6157 5843
rect -6083 5797 -6037 5843
<< polysilicon >>
rect -6960 6600 -6840 6660
rect -6720 6600 -6600 6660
rect -6480 6600 -6360 6660
rect -6240 6600 -6120 6660
rect -6960 6120 -6840 6240
rect -6720 6120 -6600 6240
rect -6480 6120 -6360 6240
rect -6240 6120 -6120 6240
rect -6960 6083 -6120 6120
rect -6960 6037 -6923 6083
rect -6877 6037 -6803 6083
rect -6757 6037 -6683 6083
rect -6637 6037 -6563 6083
rect -6517 6037 -6443 6083
rect -6397 6037 -6323 6083
rect -6277 6037 -6203 6083
rect -6157 6037 -6120 6083
rect -6960 6000 -6120 6037
rect -6960 4980 -6840 5040
rect -6720 4980 -6600 5040
rect -6480 4980 -6360 5040
rect -6240 4980 -6120 5040
rect -6960 4560 -6840 4680
rect -6720 4560 -6600 4680
rect -6960 4523 -6600 4560
rect -6960 4477 -6923 4523
rect -6877 4477 -6803 4523
rect -6757 4477 -6683 4523
rect -6637 4477 -6600 4523
rect -6960 4440 -6600 4477
rect -6480 4560 -6360 4680
rect -6240 4560 -6120 4680
rect -6480 4523 -6120 4560
rect -6480 4477 -6443 4523
rect -6397 4477 -6323 4523
rect -6277 4477 -6203 4523
rect -6157 4477 -6120 4523
rect -6480 4440 -6120 4477
rect -6960 -517 -6600 -480
rect -6960 -563 -6923 -517
rect -6877 -563 -6803 -517
rect -6757 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -600 -6600 -563
rect -6960 -720 -6840 -600
rect -6720 -720 -6600 -600
rect -6480 -517 -6120 -480
rect -6480 -563 -6443 -517
rect -6397 -563 -6323 -517
rect -6277 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -600 -6120 -563
rect -6480 -720 -6360 -600
rect -6240 -720 -6120 -600
rect -6960 -1140 -6840 -1080
rect -6720 -1140 -6600 -1080
rect -6480 -1140 -6360 -1080
rect -6240 -1140 -6120 -1080
<< polycontact >>
rect -6923 6037 -6877 6083
rect -6803 6037 -6757 6083
rect -6683 6037 -6637 6083
rect -6563 6037 -6517 6083
rect -6443 6037 -6397 6083
rect -6323 6037 -6277 6083
rect -6203 6037 -6157 6083
rect -6923 4477 -6877 4523
rect -6803 4477 -6757 4523
rect -6683 4477 -6637 4523
rect -6443 4477 -6397 4523
rect -6323 4477 -6277 4523
rect -6203 4477 -6157 4523
rect -6923 -563 -6877 -517
rect -6803 -563 -6757 -517
rect -6683 -563 -6637 -517
rect -6443 -563 -6397 -517
rect -6323 -563 -6277 -517
rect -6203 -563 -6157 -517
<< metal1 >>
rect -7200 7043 -5880 7080
rect -7200 6997 -7163 7043
rect -7117 6997 -7043 7043
rect -6997 6997 -6923 7043
rect -6877 6997 -6803 7043
rect -6757 6997 -6683 7043
rect -6637 6997 -6563 7043
rect -6517 6997 -6443 7043
rect -6397 6997 -6323 7043
rect -6277 6997 -6203 7043
rect -6157 6997 -6083 7043
rect -6037 6997 -5963 7043
rect -5917 6997 -5880 7043
rect -7200 6960 -5880 6997
rect -7200 6806 -5880 6840
rect -7200 6754 -7046 6806
rect -6994 6803 -6566 6806
rect -6514 6803 -6086 6806
rect -6994 6757 -6923 6803
rect -6877 6757 -6803 6803
rect -6757 6757 -6683 6803
rect -6637 6757 -6566 6803
rect -6514 6757 -6443 6803
rect -6397 6757 -6323 6803
rect -6277 6757 -6203 6803
rect -6157 6757 -6086 6803
rect -6994 6754 -6566 6757
rect -6514 6754 -6086 6757
rect -6034 6754 -5880 6806
rect -7200 6720 -5880 6754
rect -7080 6566 -6960 6600
rect -7080 6514 -7046 6566
rect -6994 6514 -6960 6566
rect -7080 6446 -6960 6514
rect -7080 6394 -7046 6446
rect -6994 6394 -6960 6446
rect -7080 6326 -6960 6394
rect -7080 6274 -7046 6326
rect -6994 6274 -6960 6326
rect -7080 6240 -6960 6274
rect -6840 6566 -6720 6600
rect -6840 6514 -6806 6566
rect -6754 6514 -6720 6566
rect -6840 6446 -6720 6514
rect -6840 6394 -6806 6446
rect -6754 6394 -6720 6446
rect -6840 6326 -6720 6394
rect -6840 6274 -6806 6326
rect -6754 6274 -6720 6326
rect -6840 6240 -6720 6274
rect -6600 6566 -6480 6600
rect -6600 6514 -6566 6566
rect -6514 6514 -6480 6566
rect -6600 6446 -6480 6514
rect -6600 6394 -6566 6446
rect -6514 6394 -6480 6446
rect -6600 6326 -6480 6394
rect -6600 6274 -6566 6326
rect -6514 6274 -6480 6326
rect -6600 6240 -6480 6274
rect -6360 6566 -6240 6600
rect -6360 6514 -6326 6566
rect -6274 6514 -6240 6566
rect -6360 6446 -6240 6514
rect -6360 6394 -6326 6446
rect -6274 6394 -6240 6446
rect -6360 6326 -6240 6394
rect -6360 6274 -6326 6326
rect -6274 6274 -6240 6326
rect -6360 6240 -6240 6274
rect -6120 6566 -6000 6600
rect -6120 6514 -6086 6566
rect -6034 6514 -6000 6566
rect -6120 6446 -6000 6514
rect -6120 6394 -6086 6446
rect -6034 6394 -6000 6446
rect -6120 6326 -6000 6394
rect -6120 6274 -6086 6326
rect -6034 6274 -6000 6326
rect -6120 6240 -6000 6274
rect -6960 6086 -6120 6120
rect -6960 6083 -6566 6086
rect -6514 6083 -6120 6086
rect -6960 6037 -6923 6083
rect -6877 6037 -6803 6083
rect -6757 6037 -6683 6083
rect -6637 6037 -6566 6083
rect -6514 6037 -6443 6083
rect -6397 6037 -6323 6083
rect -6277 6037 -6203 6083
rect -6157 6037 -6120 6083
rect -6960 6034 -6566 6037
rect -6514 6034 -6120 6037
rect -6960 6000 -6120 6034
rect -7200 5843 -5880 5880
rect -7200 5797 -7043 5843
rect -6997 5797 -6923 5843
rect -6877 5797 -6803 5843
rect -6757 5797 -6683 5843
rect -6637 5797 -6563 5843
rect -6517 5797 -6443 5843
rect -6397 5797 -6323 5843
rect -6277 5797 -6203 5843
rect -6157 5797 -6083 5843
rect -6037 5797 -5880 5843
rect -7200 5760 -5880 5797
rect -7200 5603 -5880 5640
rect -7200 5557 -7163 5603
rect -7117 5557 -7043 5603
rect -6997 5557 -6923 5603
rect -6877 5557 -6803 5603
rect -6757 5557 -6683 5603
rect -6637 5557 -6563 5603
rect -6517 5557 -6443 5603
rect -6397 5557 -6323 5603
rect -6277 5557 -6203 5603
rect -6157 5557 -6083 5603
rect -6037 5557 -5963 5603
rect -5917 5557 -5880 5603
rect -7200 5520 -5880 5557
rect -7200 5363 -5880 5400
rect -7200 5317 -7043 5363
rect -6997 5317 -6923 5363
rect -6877 5317 -6803 5363
rect -6757 5317 -6683 5363
rect -6637 5317 -6563 5363
rect -6517 5317 -6443 5363
rect -6397 5317 -6323 5363
rect -6277 5317 -6203 5363
rect -6157 5317 -6083 5363
rect -6037 5317 -5880 5363
rect -7200 5280 -5880 5317
rect -7080 5126 -6000 5160
rect -7080 5074 -7046 5126
rect -6994 5074 -6566 5126
rect -6514 5074 -6086 5126
rect -6034 5074 -6000 5126
rect -7080 5040 -6000 5074
rect -7080 5006 -6960 5040
rect -7080 4954 -7046 5006
rect -6994 4954 -6960 5006
rect -6600 5006 -6480 5040
rect -7080 4886 -6960 4954
rect -7080 4834 -7046 4886
rect -6994 4834 -6960 4886
rect -7080 4766 -6960 4834
rect -7080 4714 -7046 4766
rect -6994 4714 -6960 4766
rect -7080 4680 -6960 4714
rect -6840 4886 -6720 4980
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4766 -6720 4834
rect -6840 4714 -6806 4766
rect -6754 4714 -6720 4766
rect -6840 4680 -6720 4714
rect -6600 4954 -6566 5006
rect -6514 4954 -6480 5006
rect -6120 5006 -6000 5040
rect -6600 4883 -6480 4954
rect -6600 4837 -6563 4883
rect -6517 4837 -6480 4883
rect -6600 4763 -6480 4837
rect -6600 4717 -6563 4763
rect -6517 4717 -6480 4763
rect -6600 4680 -6480 4717
rect -6360 4886 -6240 4980
rect -6360 4834 -6326 4886
rect -6274 4834 -6240 4886
rect -6360 4766 -6240 4834
rect -6360 4714 -6326 4766
rect -6274 4714 -6240 4766
rect -6360 4680 -6240 4714
rect -6120 4954 -6086 5006
rect -6034 4954 -6000 5006
rect -6120 4886 -6000 4954
rect -6120 4834 -6086 4886
rect -6034 4834 -6000 4886
rect -6120 4766 -6000 4834
rect -6120 4714 -6086 4766
rect -6034 4714 -6000 4766
rect -6120 4680 -6000 4714
rect -6960 4526 -6600 4560
rect -6960 4523 -6806 4526
rect -6754 4523 -6600 4526
rect -6960 4477 -6923 4523
rect -6877 4477 -6806 4523
rect -6754 4477 -6683 4523
rect -6637 4477 -6600 4523
rect -6960 4474 -6806 4477
rect -6754 4474 -6600 4477
rect -6960 4440 -6600 4474
rect -6480 4526 -6120 4560
rect -6480 4523 -6326 4526
rect -6274 4523 -6120 4526
rect -6480 4477 -6443 4523
rect -6397 4477 -6326 4523
rect -6274 4477 -6203 4523
rect -6157 4477 -6120 4523
rect -6480 4474 -6326 4477
rect -6274 4474 -6120 4477
rect -6480 4440 -6120 4474
rect -7200 4286 -5880 4320
rect -7200 4234 -7046 4286
rect -6994 4283 -6086 4286
rect -6994 4237 -6923 4283
rect -6877 4237 -6803 4283
rect -6757 4237 -6683 4283
rect -6637 4237 -6563 4283
rect -6517 4237 -6443 4283
rect -6397 4237 -6323 4283
rect -6277 4237 -6203 4283
rect -6157 4237 -6086 4283
rect -6994 4234 -6086 4237
rect -6034 4234 -5880 4286
rect -7200 4200 -5880 4234
rect -7200 4046 -5880 4080
rect -7200 4043 -7046 4046
rect -6994 4043 -6086 4046
rect -6034 4043 -5880 4046
rect -7200 3997 -7163 4043
rect -7117 3997 -7046 4043
rect -6994 3997 -6923 4043
rect -6877 3997 -6803 4043
rect -6757 3997 -6683 4043
rect -6637 3997 -6563 4043
rect -6517 3997 -6443 4043
rect -6397 3997 -6323 4043
rect -6277 3997 -6203 4043
rect -6157 3997 -6086 4043
rect -6034 3997 -5963 4043
rect -5917 3997 -5880 4043
rect -7200 3994 -7046 3997
rect -6994 3994 -6086 3997
rect -6034 3994 -5880 3997
rect -7200 3960 -5880 3994
rect -7200 2846 -5880 2880
rect -7200 2843 -7046 2846
rect -6994 2843 -6086 2846
rect -6034 2843 -5880 2846
rect -7200 2797 -7163 2843
rect -7117 2797 -7046 2843
rect -6994 2797 -6923 2843
rect -6877 2797 -6803 2843
rect -6757 2797 -6683 2843
rect -6637 2797 -6563 2843
rect -6517 2797 -6443 2843
rect -6397 2797 -6323 2843
rect -6277 2797 -6203 2843
rect -6157 2797 -6086 2843
rect -6034 2797 -5963 2843
rect -5917 2797 -5880 2843
rect -7200 2794 -7046 2797
rect -6994 2794 -6086 2797
rect -6034 2794 -5880 2797
rect -7200 2760 -5880 2794
rect -7200 2366 -5880 2400
rect -7200 2363 -7046 2366
rect -6994 2363 -6086 2366
rect -6034 2363 -5880 2366
rect -7200 2317 -7163 2363
rect -7117 2317 -7046 2363
rect -6994 2317 -6923 2363
rect -6877 2317 -6803 2363
rect -6757 2317 -6683 2363
rect -6637 2317 -6563 2363
rect -6517 2317 -6443 2363
rect -6397 2317 -6323 2363
rect -6277 2317 -6203 2363
rect -6157 2317 -6086 2363
rect -6034 2317 -5963 2363
rect -5917 2317 -5880 2363
rect -7200 2314 -7046 2317
rect -6994 2314 -6086 2317
rect -6034 2314 -5880 2317
rect -7200 2280 -5880 2314
rect -7200 1886 -5880 1920
rect -7200 1883 -7046 1886
rect -6994 1883 -6086 1886
rect -6034 1883 -5880 1886
rect -7200 1837 -7163 1883
rect -7117 1837 -7046 1883
rect -6994 1837 -6923 1883
rect -6877 1837 -6803 1883
rect -6757 1837 -6683 1883
rect -6637 1837 -6563 1883
rect -6517 1837 -6443 1883
rect -6397 1837 -6323 1883
rect -6277 1837 -6203 1883
rect -6157 1837 -6086 1883
rect -6034 1837 -5963 1883
rect -5917 1837 -5880 1883
rect -7200 1834 -7046 1837
rect -6994 1834 -6086 1837
rect -6034 1834 -5880 1837
rect -7200 1800 -5880 1834
rect -7200 1406 -5880 1440
rect -7200 1403 -7046 1406
rect -6994 1403 -6086 1406
rect -6034 1403 -5880 1406
rect -7200 1357 -7163 1403
rect -7117 1357 -7046 1403
rect -6994 1357 -6923 1403
rect -6877 1357 -6803 1403
rect -6757 1357 -6683 1403
rect -6637 1357 -6563 1403
rect -6517 1357 -6443 1403
rect -6397 1357 -6323 1403
rect -6277 1357 -6203 1403
rect -6157 1357 -6086 1403
rect -6034 1357 -5963 1403
rect -5917 1357 -5880 1403
rect -7200 1354 -7046 1357
rect -6994 1354 -6086 1357
rect -6034 1354 -5880 1357
rect -7200 1320 -5880 1354
rect -7200 926 -5880 960
rect -7200 923 -7046 926
rect -6994 923 -6086 926
rect -6034 923 -5880 926
rect -7200 877 -7163 923
rect -7117 877 -7046 923
rect -6994 877 -6923 923
rect -6877 877 -6803 923
rect -6757 877 -6683 923
rect -6637 877 -6563 923
rect -6517 877 -6443 923
rect -6397 877 -6323 923
rect -6277 877 -6203 923
rect -6157 877 -6086 923
rect -6034 877 -5963 923
rect -5917 877 -5880 923
rect -7200 874 -7046 877
rect -6994 874 -6086 877
rect -6034 874 -5880 877
rect -7200 840 -5880 874
rect -7200 -274 -5880 -240
rect -7200 -277 -7046 -274
rect -6994 -277 -6086 -274
rect -6034 -277 -5880 -274
rect -7200 -323 -7163 -277
rect -7117 -323 -7046 -277
rect -6994 -323 -6923 -277
rect -6877 -323 -6803 -277
rect -6757 -323 -6683 -277
rect -6637 -323 -6563 -277
rect -6517 -323 -6443 -277
rect -6397 -323 -6323 -277
rect -6277 -323 -6203 -277
rect -6157 -323 -6086 -277
rect -6034 -323 -5963 -277
rect -5917 -323 -5880 -277
rect -7200 -326 -7046 -323
rect -6994 -326 -6086 -323
rect -6034 -326 -5880 -323
rect -7200 -360 -5880 -326
rect -6960 -514 -6600 -480
rect -6960 -517 -6806 -514
rect -6754 -517 -6600 -514
rect -6960 -563 -6923 -517
rect -6877 -563 -6806 -517
rect -6754 -563 -6683 -517
rect -6637 -563 -6600 -517
rect -6960 -566 -6806 -563
rect -6754 -566 -6600 -563
rect -6960 -600 -6600 -566
rect -6480 -514 -6120 -480
rect -6480 -517 -6326 -514
rect -6274 -517 -6120 -514
rect -6480 -563 -6443 -517
rect -6397 -563 -6326 -517
rect -6274 -563 -6203 -517
rect -6157 -563 -6120 -517
rect -6480 -566 -6326 -563
rect -6274 -566 -6120 -563
rect -6480 -600 -6120 -566
rect -7080 -754 -6960 -720
rect -7080 -806 -7046 -754
rect -6994 -806 -6960 -754
rect -7080 -874 -6960 -806
rect -7080 -926 -7046 -874
rect -6994 -926 -6960 -874
rect -7080 -994 -6960 -926
rect -7080 -1046 -7046 -994
rect -6994 -1046 -6960 -994
rect -7080 -1080 -6960 -1046
rect -6840 -757 -6720 -720
rect -6840 -803 -6803 -757
rect -6757 -803 -6720 -757
rect -6840 -877 -6720 -803
rect -6840 -923 -6803 -877
rect -6757 -923 -6720 -877
rect -6840 -997 -6720 -923
rect -6840 -1043 -6803 -997
rect -6757 -1043 -6720 -997
rect -6840 -1080 -6720 -1043
rect -6600 -754 -6480 -720
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6360 -757 -6240 -720
rect -6360 -803 -6323 -757
rect -6277 -803 -6240 -757
rect -6360 -877 -6240 -803
rect -6360 -923 -6323 -877
rect -6277 -923 -6240 -877
rect -6360 -997 -6240 -923
rect -6360 -1043 -6323 -997
rect -6277 -1043 -6240 -997
rect -6360 -1080 -6240 -1043
rect -6120 -754 -6000 -720
rect -6120 -806 -6086 -754
rect -6034 -806 -6000 -754
rect -6120 -874 -6000 -806
rect -6120 -926 -6086 -874
rect -6034 -926 -6000 -874
rect -6120 -994 -6000 -926
rect -6120 -1046 -6086 -994
rect -6034 -1046 -6000 -994
rect -6120 -1080 -6000 -1046
rect -7200 -1234 -5880 -1200
rect -7200 -1237 -7046 -1234
rect -6994 -1237 -6086 -1234
rect -6034 -1237 -5880 -1234
rect -7200 -1283 -7163 -1237
rect -7117 -1283 -7046 -1237
rect -6994 -1283 -6923 -1237
rect -6877 -1283 -6803 -1237
rect -6757 -1283 -6683 -1237
rect -6637 -1283 -6563 -1237
rect -6517 -1283 -6443 -1237
rect -6397 -1283 -6323 -1237
rect -6277 -1283 -6203 -1237
rect -6157 -1283 -6086 -1237
rect -6034 -1283 -5963 -1237
rect -5917 -1283 -5880 -1237
rect -7200 -1286 -7046 -1283
rect -6994 -1286 -6086 -1283
rect -6034 -1286 -5880 -1283
rect -7200 -1320 -5880 -1286
<< via1 >>
rect -7046 6803 -6994 6806
rect -6566 6803 -6514 6806
rect -6086 6803 -6034 6806
rect -7046 6757 -7043 6803
rect -7043 6757 -6997 6803
rect -6997 6757 -6994 6803
rect -6566 6757 -6563 6803
rect -6563 6757 -6517 6803
rect -6517 6757 -6514 6803
rect -6086 6757 -6083 6803
rect -6083 6757 -6037 6803
rect -6037 6757 -6034 6803
rect -7046 6754 -6994 6757
rect -6566 6754 -6514 6757
rect -6086 6754 -6034 6757
rect -7046 6563 -6994 6566
rect -7046 6517 -7043 6563
rect -7043 6517 -6997 6563
rect -6997 6517 -6994 6563
rect -7046 6514 -6994 6517
rect -7046 6443 -6994 6446
rect -7046 6397 -7043 6443
rect -7043 6397 -6997 6443
rect -6997 6397 -6994 6443
rect -7046 6394 -6994 6397
rect -7046 6323 -6994 6326
rect -7046 6277 -7043 6323
rect -7043 6277 -6997 6323
rect -6997 6277 -6994 6323
rect -7046 6274 -6994 6277
rect -6806 6563 -6754 6566
rect -6806 6517 -6803 6563
rect -6803 6517 -6757 6563
rect -6757 6517 -6754 6563
rect -6806 6514 -6754 6517
rect -6806 6443 -6754 6446
rect -6806 6397 -6803 6443
rect -6803 6397 -6757 6443
rect -6757 6397 -6754 6443
rect -6806 6394 -6754 6397
rect -6806 6323 -6754 6326
rect -6806 6277 -6803 6323
rect -6803 6277 -6757 6323
rect -6757 6277 -6754 6323
rect -6806 6274 -6754 6277
rect -6566 6563 -6514 6566
rect -6566 6517 -6563 6563
rect -6563 6517 -6517 6563
rect -6517 6517 -6514 6563
rect -6566 6514 -6514 6517
rect -6566 6443 -6514 6446
rect -6566 6397 -6563 6443
rect -6563 6397 -6517 6443
rect -6517 6397 -6514 6443
rect -6566 6394 -6514 6397
rect -6566 6323 -6514 6326
rect -6566 6277 -6563 6323
rect -6563 6277 -6517 6323
rect -6517 6277 -6514 6323
rect -6566 6274 -6514 6277
rect -6326 6563 -6274 6566
rect -6326 6517 -6323 6563
rect -6323 6517 -6277 6563
rect -6277 6517 -6274 6563
rect -6326 6514 -6274 6517
rect -6326 6443 -6274 6446
rect -6326 6397 -6323 6443
rect -6323 6397 -6277 6443
rect -6277 6397 -6274 6443
rect -6326 6394 -6274 6397
rect -6326 6323 -6274 6326
rect -6326 6277 -6323 6323
rect -6323 6277 -6277 6323
rect -6277 6277 -6274 6323
rect -6326 6274 -6274 6277
rect -6086 6563 -6034 6566
rect -6086 6517 -6083 6563
rect -6083 6517 -6037 6563
rect -6037 6517 -6034 6563
rect -6086 6514 -6034 6517
rect -6086 6443 -6034 6446
rect -6086 6397 -6083 6443
rect -6083 6397 -6037 6443
rect -6037 6397 -6034 6443
rect -6086 6394 -6034 6397
rect -6086 6323 -6034 6326
rect -6086 6277 -6083 6323
rect -6083 6277 -6037 6323
rect -6037 6277 -6034 6323
rect -6086 6274 -6034 6277
rect -6566 6083 -6514 6086
rect -6566 6037 -6563 6083
rect -6563 6037 -6517 6083
rect -6517 6037 -6514 6083
rect -6566 6034 -6514 6037
rect -7046 5074 -6994 5126
rect -6566 5074 -6514 5126
rect -6086 5074 -6034 5126
rect -7046 4954 -6994 5006
rect -7046 4883 -6994 4886
rect -7046 4837 -7043 4883
rect -7043 4837 -6997 4883
rect -6997 4837 -6994 4883
rect -7046 4834 -6994 4837
rect -7046 4763 -6994 4766
rect -7046 4717 -7043 4763
rect -7043 4717 -6997 4763
rect -6997 4717 -6994 4763
rect -7046 4714 -6994 4717
rect -6806 4883 -6754 4886
rect -6806 4837 -6803 4883
rect -6803 4837 -6757 4883
rect -6757 4837 -6754 4883
rect -6806 4834 -6754 4837
rect -6806 4763 -6754 4766
rect -6806 4717 -6803 4763
rect -6803 4717 -6757 4763
rect -6757 4717 -6754 4763
rect -6806 4714 -6754 4717
rect -6566 4954 -6514 5006
rect -6326 4883 -6274 4886
rect -6326 4837 -6323 4883
rect -6323 4837 -6277 4883
rect -6277 4837 -6274 4883
rect -6326 4834 -6274 4837
rect -6326 4763 -6274 4766
rect -6326 4717 -6323 4763
rect -6323 4717 -6277 4763
rect -6277 4717 -6274 4763
rect -6326 4714 -6274 4717
rect -6086 4954 -6034 5006
rect -6086 4883 -6034 4886
rect -6086 4837 -6083 4883
rect -6083 4837 -6037 4883
rect -6037 4837 -6034 4883
rect -6086 4834 -6034 4837
rect -6086 4763 -6034 4766
rect -6086 4717 -6083 4763
rect -6083 4717 -6037 4763
rect -6037 4717 -6034 4763
rect -6086 4714 -6034 4717
rect -6806 4523 -6754 4526
rect -6806 4477 -6803 4523
rect -6803 4477 -6757 4523
rect -6757 4477 -6754 4523
rect -6806 4474 -6754 4477
rect -6326 4523 -6274 4526
rect -6326 4477 -6323 4523
rect -6323 4477 -6277 4523
rect -6277 4477 -6274 4523
rect -6326 4474 -6274 4477
rect -7046 4283 -6994 4286
rect -6086 4283 -6034 4286
rect -7046 4237 -7043 4283
rect -7043 4237 -6997 4283
rect -6997 4237 -6994 4283
rect -6086 4237 -6083 4283
rect -6083 4237 -6037 4283
rect -6037 4237 -6034 4283
rect -7046 4234 -6994 4237
rect -6086 4234 -6034 4237
rect -7046 4043 -6994 4046
rect -6086 4043 -6034 4046
rect -7046 3997 -7043 4043
rect -7043 3997 -6997 4043
rect -6997 3997 -6994 4043
rect -6086 3997 -6083 4043
rect -6083 3997 -6037 4043
rect -6037 3997 -6034 4043
rect -7046 3994 -6994 3997
rect -6086 3994 -6034 3997
rect -7046 2843 -6994 2846
rect -6086 2843 -6034 2846
rect -7046 2797 -7043 2843
rect -7043 2797 -6997 2843
rect -6997 2797 -6994 2843
rect -6086 2797 -6083 2843
rect -6083 2797 -6037 2843
rect -6037 2797 -6034 2843
rect -7046 2794 -6994 2797
rect -6086 2794 -6034 2797
rect -7046 2363 -6994 2366
rect -6086 2363 -6034 2366
rect -7046 2317 -7043 2363
rect -7043 2317 -6997 2363
rect -6997 2317 -6994 2363
rect -6086 2317 -6083 2363
rect -6083 2317 -6037 2363
rect -6037 2317 -6034 2363
rect -7046 2314 -6994 2317
rect -6086 2314 -6034 2317
rect -7046 1883 -6994 1886
rect -6086 1883 -6034 1886
rect -7046 1837 -7043 1883
rect -7043 1837 -6997 1883
rect -6997 1837 -6994 1883
rect -6086 1837 -6083 1883
rect -6083 1837 -6037 1883
rect -6037 1837 -6034 1883
rect -7046 1834 -6994 1837
rect -6086 1834 -6034 1837
rect -7046 1403 -6994 1406
rect -6086 1403 -6034 1406
rect -7046 1357 -7043 1403
rect -7043 1357 -6997 1403
rect -6997 1357 -6994 1403
rect -6086 1357 -6083 1403
rect -6083 1357 -6037 1403
rect -6037 1357 -6034 1403
rect -7046 1354 -6994 1357
rect -6086 1354 -6034 1357
rect -7046 923 -6994 926
rect -6086 923 -6034 926
rect -7046 877 -7043 923
rect -7043 877 -6997 923
rect -6997 877 -6994 923
rect -6086 877 -6083 923
rect -6083 877 -6037 923
rect -6037 877 -6034 923
rect -7046 874 -6994 877
rect -6086 874 -6034 877
rect -7046 -277 -6994 -274
rect -6086 -277 -6034 -274
rect -7046 -323 -7043 -277
rect -7043 -323 -6997 -277
rect -6997 -323 -6994 -277
rect -6086 -323 -6083 -277
rect -6083 -323 -6037 -277
rect -6037 -323 -6034 -277
rect -7046 -326 -6994 -323
rect -6086 -326 -6034 -323
rect -6806 -517 -6754 -514
rect -6806 -563 -6803 -517
rect -6803 -563 -6757 -517
rect -6757 -563 -6754 -517
rect -6806 -566 -6754 -563
rect -6326 -517 -6274 -514
rect -6326 -563 -6323 -517
rect -6323 -563 -6277 -517
rect -6277 -563 -6274 -517
rect -6326 -566 -6274 -563
rect -7046 -757 -6994 -754
rect -7046 -803 -7043 -757
rect -7043 -803 -6997 -757
rect -6997 -803 -6994 -757
rect -7046 -806 -6994 -803
rect -7046 -877 -6994 -874
rect -7046 -923 -7043 -877
rect -7043 -923 -6997 -877
rect -6997 -923 -6994 -877
rect -7046 -926 -6994 -923
rect -7046 -997 -6994 -994
rect -7046 -1043 -7043 -997
rect -7043 -1043 -6997 -997
rect -6997 -1043 -6994 -997
rect -7046 -1046 -6994 -1043
rect -6566 -757 -6514 -754
rect -6566 -803 -6563 -757
rect -6563 -803 -6517 -757
rect -6517 -803 -6514 -757
rect -6566 -806 -6514 -803
rect -6566 -877 -6514 -874
rect -6566 -923 -6563 -877
rect -6563 -923 -6517 -877
rect -6517 -923 -6514 -877
rect -6566 -926 -6514 -923
rect -6566 -997 -6514 -994
rect -6566 -1043 -6563 -997
rect -6563 -1043 -6517 -997
rect -6517 -1043 -6514 -997
rect -6566 -1046 -6514 -1043
rect -6086 -757 -6034 -754
rect -6086 -803 -6083 -757
rect -6083 -803 -6037 -757
rect -6037 -803 -6034 -757
rect -6086 -806 -6034 -803
rect -6086 -877 -6034 -874
rect -6086 -923 -6083 -877
rect -6083 -923 -6037 -877
rect -6037 -923 -6034 -877
rect -6086 -926 -6034 -923
rect -6086 -997 -6034 -994
rect -6086 -1043 -6083 -997
rect -6083 -1043 -6037 -997
rect -6037 -1043 -6034 -997
rect -6086 -1046 -6034 -1043
rect -7046 -1237 -6994 -1234
rect -6086 -1237 -6034 -1234
rect -7046 -1283 -7043 -1237
rect -7043 -1283 -6997 -1237
rect -6997 -1283 -6994 -1237
rect -6086 -1283 -6083 -1237
rect -6083 -1283 -6037 -1237
rect -6037 -1283 -6034 -1237
rect -7046 -1286 -6994 -1283
rect -6086 -1286 -6034 -1283
<< metal2 >>
rect -7080 6808 -6960 6840
rect -7080 6752 -7048 6808
rect -6992 6752 -6960 6808
rect -7080 6568 -6960 6752
rect -6600 6808 -6480 6840
rect -6600 6752 -6568 6808
rect -6512 6752 -6480 6808
rect -7080 6512 -7048 6568
rect -6992 6512 -6960 6568
rect -7080 6448 -6960 6512
rect -7080 6392 -7048 6448
rect -6992 6392 -6960 6448
rect -7080 6328 -6960 6392
rect -7080 6272 -7048 6328
rect -6992 6272 -6960 6328
rect -7080 6240 -6960 6272
rect -6840 6566 -6720 6600
rect -6840 6514 -6806 6566
rect -6754 6514 -6720 6566
rect -6840 6446 -6720 6514
rect -6840 6394 -6806 6446
rect -6754 6394 -6720 6446
rect -6840 6326 -6720 6394
rect -6840 6274 -6806 6326
rect -6754 6274 -6720 6326
rect -6840 5848 -6720 6274
rect -6600 6568 -6480 6752
rect -6120 6808 -6000 6840
rect -6120 6752 -6088 6808
rect -6032 6752 -6000 6808
rect -6600 6512 -6568 6568
rect -6512 6512 -6480 6568
rect -6600 6448 -6480 6512
rect -6600 6392 -6568 6448
rect -6512 6392 -6480 6448
rect -6600 6328 -6480 6392
rect -6600 6272 -6568 6328
rect -6512 6272 -6480 6328
rect -6600 6240 -6480 6272
rect -6360 6566 -6240 6600
rect -6360 6514 -6326 6566
rect -6274 6514 -6240 6566
rect -6360 6446 -6240 6514
rect -6360 6394 -6326 6446
rect -6274 6394 -6240 6446
rect -6360 6326 -6240 6394
rect -6360 6274 -6326 6326
rect -6274 6274 -6240 6326
rect -6600 6088 -6480 6120
rect -6600 6032 -6568 6088
rect -6512 6032 -6480 6088
rect -6600 6000 -6480 6032
rect -6840 5792 -6808 5848
rect -6752 5792 -6720 5848
rect -7080 5368 -6960 5400
rect -7080 5312 -7048 5368
rect -6992 5312 -6960 5368
rect -7080 5126 -6960 5312
rect -6840 5368 -6720 5792
rect -6360 5848 -6240 6274
rect -6120 6568 -6000 6752
rect -6120 6512 -6088 6568
rect -6032 6512 -6000 6568
rect -6120 6448 -6000 6512
rect -6120 6392 -6088 6448
rect -6032 6392 -6000 6448
rect -6120 6328 -6000 6392
rect -6120 6272 -6088 6328
rect -6032 6272 -6000 6328
rect -6120 6240 -6000 6272
rect -6360 5792 -6328 5848
rect -6272 5792 -6240 5848
rect -6840 5312 -6808 5368
rect -6752 5312 -6720 5368
rect -6840 5280 -6720 5312
rect -6600 5368 -6480 5400
rect -6600 5312 -6568 5368
rect -6512 5312 -6480 5368
rect -7080 5074 -7046 5126
rect -6994 5074 -6960 5126
rect -7080 5006 -6960 5074
rect -7080 4954 -7046 5006
rect -6994 4954 -6960 5006
rect -6600 5126 -6480 5312
rect -6360 5368 -6240 5792
rect -6360 5312 -6328 5368
rect -6272 5312 -6240 5368
rect -6360 5280 -6240 5312
rect -6120 5368 -6000 5400
rect -6120 5312 -6088 5368
rect -6032 5312 -6000 5368
rect -6600 5074 -6566 5126
rect -6514 5074 -6480 5126
rect -6600 5006 -6480 5074
rect -7080 4886 -6960 4954
rect -7080 4834 -7046 4886
rect -6994 4834 -6960 4886
rect -7080 4766 -6960 4834
rect -7080 4714 -7046 4766
rect -6994 4714 -6960 4766
rect -7080 4680 -6960 4714
rect -6840 4886 -6720 4980
rect -6600 4954 -6566 5006
rect -6514 4954 -6480 5006
rect -6120 5126 -6000 5312
rect -6120 5074 -6086 5126
rect -6034 5074 -6000 5126
rect -6120 5006 -6000 5074
rect -6600 4920 -6480 4954
rect -6840 4834 -6806 4886
rect -6754 4834 -6720 4886
rect -6840 4800 -6720 4834
rect -6360 4886 -6240 4980
rect -6360 4834 -6326 4886
rect -6274 4834 -6240 4886
rect -6360 4800 -6240 4834
rect -6840 4766 -6240 4800
rect -6840 4714 -6806 4766
rect -6754 4714 -6326 4766
rect -6274 4714 -6240 4766
rect -6840 4680 -6240 4714
rect -6120 4954 -6086 5006
rect -6034 4954 -6000 5006
rect -6120 4886 -6000 4954
rect -6120 4834 -6086 4886
rect -6034 4834 -6000 4886
rect -6120 4766 -6000 4834
rect -6120 4714 -6086 4766
rect -6034 4714 -6000 4766
rect -6120 4680 -6000 4714
rect -6840 4528 -6720 4560
rect -6840 4472 -6808 4528
rect -6752 4472 -6720 4528
rect -6840 4440 -6720 4472
rect -7080 4288 -6960 4320
rect -7080 4232 -7048 4288
rect -6992 4232 -6960 4288
rect -7080 4200 -6960 4232
rect -7080 4048 -6960 4080
rect -7080 3992 -7048 4048
rect -6992 3992 -6960 4048
rect -7080 2848 -6960 3992
rect -7080 2792 -7048 2848
rect -6992 2792 -6960 2848
rect -7080 2368 -6960 2792
rect -7080 2312 -7048 2368
rect -6992 2312 -6960 2368
rect -7080 1888 -6960 2312
rect -7080 1832 -7048 1888
rect -6992 1832 -6960 1888
rect -7080 1408 -6960 1832
rect -7080 1352 -7048 1408
rect -6992 1352 -6960 1408
rect -7080 928 -6960 1352
rect -7080 872 -7048 928
rect -6992 872 -6960 928
rect -7080 -272 -6960 872
rect -7080 -328 -7048 -272
rect -6992 -328 -6960 -272
rect -7080 -752 -6960 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -7080 -808 -7048 -752
rect -6992 -808 -6960 -752
rect -7080 -872 -6960 -808
rect -7080 -928 -7048 -872
rect -6992 -928 -6960 -872
rect -7080 -992 -6960 -928
rect -7080 -1048 -7048 -992
rect -6992 -1048 -6960 -992
rect -7080 -1232 -6960 -1048
rect -6600 -754 -6480 4680
rect -6360 4528 -6240 4560
rect -6360 4472 -6328 4528
rect -6272 4472 -6240 4528
rect -6360 4440 -6240 4472
rect -6120 4288 -6000 4320
rect -6120 4232 -6088 4288
rect -6032 4232 -6000 4288
rect -6120 4200 -6000 4232
rect -6120 4048 -6000 4080
rect -6120 3992 -6088 4048
rect -6032 3992 -6000 4048
rect -6120 2848 -6000 3992
rect -6120 2792 -6088 2848
rect -6032 2792 -6000 2848
rect -6120 2368 -6000 2792
rect -6120 2312 -6088 2368
rect -6032 2312 -6000 2368
rect -6120 1888 -6000 2312
rect -6120 1832 -6088 1888
rect -6032 1832 -6000 1888
rect -6120 1408 -6000 1832
rect -6120 1352 -6088 1408
rect -6032 1352 -6000 1408
rect -6120 928 -6000 1352
rect -6120 872 -6088 928
rect -6032 872 -6000 928
rect -6120 -272 -6000 872
rect -6120 -328 -6088 -272
rect -6032 -328 -6000 -272
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -6600 -806 -6566 -754
rect -6514 -806 -6480 -754
rect -6600 -874 -6480 -806
rect -6600 -926 -6566 -874
rect -6514 -926 -6480 -874
rect -6600 -994 -6480 -926
rect -6600 -1046 -6566 -994
rect -6514 -1046 -6480 -994
rect -6600 -1080 -6480 -1046
rect -6120 -752 -6000 -328
rect -6120 -808 -6088 -752
rect -6032 -808 -6000 -752
rect -6120 -872 -6000 -808
rect -6120 -928 -6088 -872
rect -6032 -928 -6000 -872
rect -6120 -992 -6000 -928
rect -6120 -1048 -6088 -992
rect -6032 -1048 -6000 -992
rect -7080 -1288 -7048 -1232
rect -6992 -1288 -6960 -1232
rect -7080 -1320 -6960 -1288
rect -6120 -1232 -6000 -1048
rect -6120 -1288 -6088 -1232
rect -6032 -1288 -6000 -1232
rect -6120 -1320 -6000 -1288
<< via2 >>
rect -7048 6806 -6992 6808
rect -7048 6754 -7046 6806
rect -7046 6754 -6994 6806
rect -6994 6754 -6992 6806
rect -7048 6752 -6992 6754
rect -6568 6806 -6512 6808
rect -6568 6754 -6566 6806
rect -6566 6754 -6514 6806
rect -6514 6754 -6512 6806
rect -6568 6752 -6512 6754
rect -7048 6566 -6992 6568
rect -7048 6514 -7046 6566
rect -7046 6514 -6994 6566
rect -6994 6514 -6992 6566
rect -7048 6512 -6992 6514
rect -7048 6446 -6992 6448
rect -7048 6394 -7046 6446
rect -7046 6394 -6994 6446
rect -6994 6394 -6992 6446
rect -7048 6392 -6992 6394
rect -7048 6326 -6992 6328
rect -7048 6274 -7046 6326
rect -7046 6274 -6994 6326
rect -6994 6274 -6992 6326
rect -7048 6272 -6992 6274
rect -6088 6806 -6032 6808
rect -6088 6754 -6086 6806
rect -6086 6754 -6034 6806
rect -6034 6754 -6032 6806
rect -6088 6752 -6032 6754
rect -6568 6566 -6512 6568
rect -6568 6514 -6566 6566
rect -6566 6514 -6514 6566
rect -6514 6514 -6512 6566
rect -6568 6512 -6512 6514
rect -6568 6446 -6512 6448
rect -6568 6394 -6566 6446
rect -6566 6394 -6514 6446
rect -6514 6394 -6512 6446
rect -6568 6392 -6512 6394
rect -6568 6326 -6512 6328
rect -6568 6274 -6566 6326
rect -6566 6274 -6514 6326
rect -6514 6274 -6512 6326
rect -6568 6272 -6512 6274
rect -6568 6086 -6512 6088
rect -6568 6034 -6566 6086
rect -6566 6034 -6514 6086
rect -6514 6034 -6512 6086
rect -6568 6032 -6512 6034
rect -6808 5792 -6752 5848
rect -7048 5312 -6992 5368
rect -6088 6566 -6032 6568
rect -6088 6514 -6086 6566
rect -6086 6514 -6034 6566
rect -6034 6514 -6032 6566
rect -6088 6512 -6032 6514
rect -6088 6446 -6032 6448
rect -6088 6394 -6086 6446
rect -6086 6394 -6034 6446
rect -6034 6394 -6032 6446
rect -6088 6392 -6032 6394
rect -6088 6326 -6032 6328
rect -6088 6274 -6086 6326
rect -6086 6274 -6034 6326
rect -6034 6274 -6032 6326
rect -6088 6272 -6032 6274
rect -6328 5792 -6272 5848
rect -6808 5312 -6752 5368
rect -6568 5312 -6512 5368
rect -6328 5312 -6272 5368
rect -6088 5312 -6032 5368
rect -6808 4526 -6752 4528
rect -6808 4474 -6806 4526
rect -6806 4474 -6754 4526
rect -6754 4474 -6752 4526
rect -6808 4472 -6752 4474
rect -7048 4286 -6992 4288
rect -7048 4234 -7046 4286
rect -7046 4234 -6994 4286
rect -6994 4234 -6992 4286
rect -7048 4232 -6992 4234
rect -7048 4046 -6992 4048
rect -7048 3994 -7046 4046
rect -7046 3994 -6994 4046
rect -6994 3994 -6992 4046
rect -7048 3992 -6992 3994
rect -7048 2846 -6992 2848
rect -7048 2794 -7046 2846
rect -7046 2794 -6994 2846
rect -6994 2794 -6992 2846
rect -7048 2792 -6992 2794
rect -7048 2366 -6992 2368
rect -7048 2314 -7046 2366
rect -7046 2314 -6994 2366
rect -6994 2314 -6992 2366
rect -7048 2312 -6992 2314
rect -7048 1886 -6992 1888
rect -7048 1834 -7046 1886
rect -7046 1834 -6994 1886
rect -6994 1834 -6992 1886
rect -7048 1832 -6992 1834
rect -7048 1406 -6992 1408
rect -7048 1354 -7046 1406
rect -7046 1354 -6994 1406
rect -6994 1354 -6992 1406
rect -7048 1352 -6992 1354
rect -7048 926 -6992 928
rect -7048 874 -7046 926
rect -7046 874 -6994 926
rect -6994 874 -6992 926
rect -7048 872 -6992 874
rect -7048 -274 -6992 -272
rect -7048 -326 -7046 -274
rect -7046 -326 -6994 -274
rect -6994 -326 -6992 -274
rect -7048 -328 -6992 -326
rect -6808 -514 -6752 -512
rect -6808 -566 -6806 -514
rect -6806 -566 -6754 -514
rect -6754 -566 -6752 -514
rect -6808 -568 -6752 -566
rect -7048 -754 -6992 -752
rect -7048 -806 -7046 -754
rect -7046 -806 -6994 -754
rect -6994 -806 -6992 -754
rect -7048 -808 -6992 -806
rect -7048 -874 -6992 -872
rect -7048 -926 -7046 -874
rect -7046 -926 -6994 -874
rect -6994 -926 -6992 -874
rect -7048 -928 -6992 -926
rect -7048 -994 -6992 -992
rect -7048 -1046 -7046 -994
rect -7046 -1046 -6994 -994
rect -6994 -1046 -6992 -994
rect -7048 -1048 -6992 -1046
rect -6328 4526 -6272 4528
rect -6328 4474 -6326 4526
rect -6326 4474 -6274 4526
rect -6274 4474 -6272 4526
rect -6328 4472 -6272 4474
rect -6088 4286 -6032 4288
rect -6088 4234 -6086 4286
rect -6086 4234 -6034 4286
rect -6034 4234 -6032 4286
rect -6088 4232 -6032 4234
rect -6088 4046 -6032 4048
rect -6088 3994 -6086 4046
rect -6086 3994 -6034 4046
rect -6034 3994 -6032 4046
rect -6088 3992 -6032 3994
rect -6088 2846 -6032 2848
rect -6088 2794 -6086 2846
rect -6086 2794 -6034 2846
rect -6034 2794 -6032 2846
rect -6088 2792 -6032 2794
rect -6088 2366 -6032 2368
rect -6088 2314 -6086 2366
rect -6086 2314 -6034 2366
rect -6034 2314 -6032 2366
rect -6088 2312 -6032 2314
rect -6088 1886 -6032 1888
rect -6088 1834 -6086 1886
rect -6086 1834 -6034 1886
rect -6034 1834 -6032 1886
rect -6088 1832 -6032 1834
rect -6088 1406 -6032 1408
rect -6088 1354 -6086 1406
rect -6086 1354 -6034 1406
rect -6034 1354 -6032 1406
rect -6088 1352 -6032 1354
rect -6088 926 -6032 928
rect -6088 874 -6086 926
rect -6086 874 -6034 926
rect -6034 874 -6032 926
rect -6088 872 -6032 874
rect -6088 -274 -6032 -272
rect -6088 -326 -6086 -274
rect -6086 -326 -6034 -274
rect -6034 -326 -6032 -274
rect -6088 -328 -6032 -326
rect -6328 -514 -6272 -512
rect -6328 -566 -6326 -514
rect -6326 -566 -6274 -514
rect -6274 -566 -6272 -514
rect -6328 -568 -6272 -566
rect -6088 -754 -6032 -752
rect -6088 -806 -6086 -754
rect -6086 -806 -6034 -754
rect -6034 -806 -6032 -754
rect -6088 -808 -6032 -806
rect -6088 -874 -6032 -872
rect -6088 -926 -6086 -874
rect -6086 -926 -6034 -874
rect -6034 -926 -6032 -874
rect -6088 -928 -6032 -926
rect -6088 -994 -6032 -992
rect -6088 -1046 -6086 -994
rect -6086 -1046 -6034 -994
rect -6034 -1046 -6032 -994
rect -6088 -1048 -6032 -1046
rect -7048 -1234 -6992 -1232
rect -7048 -1286 -7046 -1234
rect -7046 -1286 -6994 -1234
rect -6994 -1286 -6992 -1234
rect -7048 -1288 -6992 -1286
rect -6088 -1234 -6032 -1232
rect -6088 -1286 -6086 -1234
rect -6086 -1286 -6034 -1234
rect -6034 -1286 -6032 -1234
rect -6088 -1288 -6032 -1286
<< metal3 >>
rect -7200 6808 -5880 6840
rect -7200 6752 -7048 6808
rect -6992 6752 -6568 6808
rect -6512 6752 -6088 6808
rect -6032 6752 -5880 6808
rect -7200 6568 -5880 6752
rect -7200 6512 -7048 6568
rect -6992 6512 -6568 6568
rect -6512 6512 -6088 6568
rect -6032 6512 -5880 6568
rect -7200 6448 -5880 6512
rect -7200 6392 -7048 6448
rect -6992 6392 -6568 6448
rect -6512 6392 -6088 6448
rect -6032 6392 -5880 6448
rect -7200 6328 -5880 6392
rect -7200 6272 -7048 6328
rect -6992 6272 -6568 6328
rect -6512 6272 -6088 6328
rect -6032 6272 -5880 6328
rect -7200 6240 -5880 6272
rect -6600 6088 -6480 6120
rect -6600 6032 -6568 6088
rect -6512 6032 -6480 6088
rect -6600 6000 -6480 6032
rect -7200 5848 -5880 5880
rect -7200 5792 -6808 5848
rect -6752 5792 -6328 5848
rect -6272 5792 -5880 5848
rect -7200 5700 -5880 5792
rect -7200 5608 -5880 5640
rect -7200 5552 -6568 5608
rect -6512 5552 -5880 5608
rect -7200 5520 -5880 5552
rect -7200 5368 -5880 5460
rect -7200 5312 -7048 5368
rect -6992 5312 -6808 5368
rect -6752 5312 -6568 5368
rect -6512 5312 -6328 5368
rect -6272 5312 -6088 5368
rect -6032 5312 -5880 5368
rect -7200 5280 -5880 5312
rect -6840 4528 -6720 4560
rect -6840 4472 -6808 4528
rect -6752 4472 -6720 4528
rect -6840 4440 -6720 4472
rect -6360 4528 -6240 4560
rect -6360 4472 -6328 4528
rect -6272 4472 -6240 4528
rect -6360 4440 -6240 4472
rect -7200 4288 -5880 4320
rect -7200 4232 -7048 4288
rect -6992 4232 -6088 4288
rect -6032 4232 -5880 4288
rect -7200 4200 -5880 4232
rect -7200 4048 -5880 4080
rect -7200 3992 -7048 4048
rect -6992 3992 -6088 4048
rect -6032 3992 -5880 4048
rect -7200 3960 -5880 3992
rect -7200 3540 -5880 3840
rect -7200 3360 -5880 3480
rect -7200 3000 -5880 3300
rect -7200 2848 -5880 2880
rect -7200 2792 -7048 2848
rect -6992 2792 -6088 2848
rect -6032 2792 -5880 2848
rect -7200 2760 -5880 2792
rect -7200 2520 -5880 2640
rect -7200 2368 -5880 2400
rect -7200 2312 -7048 2368
rect -6992 2312 -6088 2368
rect -6032 2312 -5880 2368
rect -7200 2280 -5880 2312
rect -7200 2040 -5880 2160
rect -7200 1888 -5880 1920
rect -7200 1832 -7048 1888
rect -6992 1832 -6088 1888
rect -6032 1832 -5880 1888
rect -7200 1800 -5880 1832
rect -7200 1560 -5880 1680
rect -7200 1408 -5880 1440
rect -7200 1352 -7048 1408
rect -6992 1352 -6088 1408
rect -6032 1352 -5880 1408
rect -7200 1320 -5880 1352
rect -7200 1080 -5880 1200
rect -7200 928 -5880 960
rect -7200 872 -7048 928
rect -6992 872 -6088 928
rect -6032 872 -5880 928
rect -7200 840 -5880 872
rect -7200 420 -5880 720
rect -7200 240 -5880 360
rect -7200 -120 -5880 180
rect -7200 -272 -5880 -240
rect -7200 -328 -7048 -272
rect -6992 -328 -6088 -272
rect -6032 -328 -5880 -272
rect -7200 -360 -5880 -328
rect -6840 -512 -6720 -480
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 -512 -6240 -480
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
rect -7200 -752 -5880 -720
rect -7200 -808 -7048 -752
rect -6992 -808 -6088 -752
rect -6032 -808 -5880 -752
rect -7200 -872 -5880 -808
rect -7200 -928 -7048 -872
rect -6992 -928 -6088 -872
rect -6032 -928 -5880 -872
rect -7200 -992 -5880 -928
rect -7200 -1048 -7048 -992
rect -6992 -1048 -6088 -992
rect -6032 -1048 -5880 -992
rect -7200 -1232 -5880 -1048
rect -7200 -1288 -7048 -1232
rect -6992 -1288 -6088 -1232
rect -6032 -1288 -5880 -1232
rect -7200 -1320 -5880 -1288
<< via3 >>
rect -6568 6032 -6512 6088
rect -6808 5792 -6752 5848
rect -6328 5792 -6272 5848
rect -6568 5552 -6512 5608
rect -7048 5312 -6992 5368
rect -6808 5312 -6752 5368
rect -6328 5312 -6272 5368
rect -6088 5312 -6032 5368
rect -6808 4472 -6752 4528
rect -6328 4472 -6272 4528
rect -6808 -568 -6752 -512
rect -6328 -568 -6272 -512
<< metal4 >>
rect -6600 6088 -6480 6120
rect -6600 6032 -6568 6088
rect -6512 6032 -6480 6088
rect -6840 5848 -6720 5880
rect -6840 5792 -6808 5848
rect -6752 5792 -6720 5848
rect -7080 5368 -6960 5400
rect -7080 5312 -7048 5368
rect -6992 5312 -6960 5368
rect -7080 5280 -6960 5312
rect -6840 5368 -6720 5792
rect -6600 5608 -6480 6032
rect -6600 5552 -6568 5608
rect -6512 5552 -6480 5608
rect -6600 5520 -6480 5552
rect -6360 5848 -6240 5880
rect -6360 5792 -6328 5848
rect -6272 5792 -6240 5848
rect -6840 5312 -6808 5368
rect -6752 5312 -6720 5368
rect -6840 5280 -6720 5312
rect -6360 5368 -6240 5792
rect -6360 5312 -6328 5368
rect -6272 5312 -6240 5368
rect -6360 5280 -6240 5312
rect -6120 5368 -6000 5400
rect -6120 5312 -6088 5368
rect -6032 5312 -6000 5368
rect -6120 5280 -6000 5312
rect -6840 4528 -6720 4560
rect -6840 4472 -6808 4528
rect -6752 4472 -6720 4528
rect -6840 4320 -6720 4472
rect -7080 4200 -6720 4320
rect -6840 -512 -6720 4200
rect -6840 -568 -6808 -512
rect -6752 -568 -6720 -512
rect -6840 -600 -6720 -568
rect -6360 4528 -6240 4560
rect -6360 4472 -6328 4528
rect -6272 4472 -6240 4528
rect -6360 4320 -6240 4472
rect -6360 4200 -6000 4320
rect -6360 -512 -6240 4200
rect -6360 -568 -6328 -512
rect -6272 -568 -6240 -512
rect -6360 -600 -6240 -568
<< labels >>
rlabel metal1 s -6780 -900 -6780 -900 4 dl
rlabel metal1 s -6300 -900 -6300 -900 4 dr
rlabel metal1 s -7020 5580 -7020 5580 4 gnd
rlabel metal1 s -7020 7020 -7020 7020 4 gnd
rlabel metal4 s -6840 -120 -6720 2400 4 inl
port 1 nsew
rlabel metal4 s -6360 -120 -6240 2400 4 inr
port 2 nsew
rlabel metal2 s -6600 -120 -6480 2400 4 out
port 3 nsew
rlabel metal3 s -7200 6240 -5880 6840 4 vdd
port 4 nsew
rlabel metal3 s -7200 5520 -7080 5640 4 gp
port 5 nsew
rlabel metal3 s -7200 4200 -7080 4320 4 bp
port 6 nsew
rlabel metal3 s -7200 5760 -7080 5880 4 vreg
port 7 nsew
rlabel metal3 s -7200 3720 -5880 3840 4 op
port 8 nsew
rlabel metal3 s -7200 3000 -5880 3120 4 op
port 8 nsew
rlabel metal3 s -7200 3360 -5880 3480 4 xm
port 9 nsew
rlabel metal3 s -7200 2520 -5880 2640 4 im
port 10 nsew
rlabel metal3 s -7200 1080 -5880 1200 4 ip
port 11 nsew
rlabel metal3 s -7200 240 -5880 360 4 xp
port 12 nsew
rlabel metal3 s -7200 -1320 -5880 -720 4 gnd
port 13 nsew
rlabel metal3 s -7200 -120 -5880 0 4 om
port 14 nsew
rlabel metal3 s -7200 600 -5880 720 4 om
port 14 nsew
rlabel metal3 s -7200 2040 -5880 2160 4 x
port 15 nsew
rlabel metal3 s -7200 1560 -5880 1680 4 y
port 16 nsew
<< end >>
