magic
tech gf180mcuC
magscale 1 5
timestamp 1665299846
<< error_p >>
rect 25908 8332 25992 8352
rect 25908 8324 25928 8332
rect 25936 8324 25964 8332
rect 25972 8324 25992 8332
rect 26028 8332 26112 8352
rect 26028 8324 26048 8332
rect 26056 8324 26084 8332
rect 26092 8324 26112 8332
rect 26148 8332 26232 8352
rect 26148 8324 26168 8332
rect 26176 8324 26204 8332
rect 26212 8324 26232 8332
rect 26268 8332 26352 8352
rect 26268 8324 26288 8332
rect 26296 8324 26324 8332
rect 26332 8324 26352 8332
rect 26388 8332 26472 8352
rect 26388 8324 26408 8332
rect 26416 8324 26444 8332
rect 26452 8324 26472 8332
rect 26508 8332 26592 8352
rect 26508 8324 26528 8332
rect 26536 8324 26564 8332
rect 26572 8324 26592 8332
rect 26628 8332 26712 8352
rect 26628 8324 26648 8332
rect 26656 8324 26684 8332
rect 26692 8324 26712 8332
rect 26748 8332 26832 8352
rect 26748 8324 26768 8332
rect 26776 8324 26804 8332
rect 26812 8324 26832 8332
rect 26868 8332 26952 8352
rect 26868 8324 26888 8332
rect 26896 8324 26924 8332
rect 26932 8324 26952 8332
rect 26988 8332 27072 8352
rect 26988 8324 27008 8332
rect 27016 8324 27044 8332
rect 27052 8324 27072 8332
rect 27108 8332 27192 8352
rect 27108 8324 27128 8332
rect 27136 8324 27164 8332
rect 27172 8324 27192 8332
rect 27228 8332 27312 8352
rect 27228 8324 27248 8332
rect 27256 8324 27284 8332
rect 27292 8324 27312 8332
rect 27348 8332 27432 8352
rect 27348 8324 27368 8332
rect 27376 8324 27404 8332
rect 27412 8324 27432 8332
rect 27468 8332 27552 8352
rect 27468 8324 27488 8332
rect 27496 8324 27524 8332
rect 27532 8324 27552 8332
rect 27588 8332 27672 8352
rect 27588 8324 27608 8332
rect 27616 8324 27644 8332
rect 27652 8324 27672 8332
rect 27708 8332 27792 8352
rect 27708 8324 27728 8332
rect 27736 8324 27764 8332
rect 27772 8324 27792 8332
rect 27828 8332 27912 8352
rect 27828 8324 27848 8332
rect 27856 8324 27884 8332
rect 27892 8324 27912 8332
rect 27948 8332 28032 8352
rect 27948 8324 27968 8332
rect 27976 8324 28004 8332
rect 28012 8324 28032 8332
rect 28068 8332 28152 8352
rect 28068 8324 28088 8332
rect 28096 8324 28124 8332
rect 28132 8324 28152 8332
rect 28188 8332 28272 8352
rect 28188 8324 28208 8332
rect 28216 8324 28244 8332
rect 28252 8324 28272 8332
rect 28308 8332 28392 8352
rect 28308 8324 28328 8332
rect 28336 8324 28364 8332
rect 28372 8324 28392 8332
rect 28428 8332 28512 8352
rect 28428 8324 28448 8332
rect 28456 8324 28484 8332
rect 28492 8324 28512 8332
rect 28548 8332 28632 8352
rect 28548 8324 28568 8332
rect 28576 8324 28604 8332
rect 28612 8324 28632 8332
rect 28668 8332 28752 8352
rect 28668 8324 28688 8332
rect 28696 8324 28724 8332
rect 28732 8324 28752 8332
rect 28788 8332 28872 8352
rect 28788 8324 28808 8332
rect 28816 8324 28844 8332
rect 28852 8324 28872 8332
rect 28908 8332 28992 8352
rect 28908 8324 28928 8332
rect 28936 8324 28964 8332
rect 28972 8324 28992 8332
rect 29028 8332 29112 8352
rect 29028 8324 29048 8332
rect 29056 8324 29084 8332
rect 29092 8324 29112 8332
rect 29148 8332 29232 8352
rect 29148 8324 29168 8332
rect 29176 8324 29204 8332
rect 29212 8324 29232 8332
rect 29268 8332 29352 8352
rect 29268 8324 29288 8332
rect 29296 8324 29324 8332
rect 29332 8324 29352 8332
rect 29388 8332 29472 8352
rect 29388 8324 29408 8332
rect 29416 8324 29444 8332
rect 29452 8324 29472 8332
rect 29508 8332 29592 8352
rect 29508 8324 29528 8332
rect 29536 8324 29564 8332
rect 29572 8324 29592 8332
rect 29628 8332 29712 8352
rect 29628 8324 29648 8332
rect 29656 8324 29684 8332
rect 29692 8324 29712 8332
rect 29748 8332 29832 8352
rect 29748 8324 29768 8332
rect 29776 8324 29804 8332
rect 29812 8324 29832 8332
rect 29868 8332 29952 8352
rect 29868 8324 29888 8332
rect 29896 8324 29924 8332
rect 29932 8324 29952 8332
rect 29988 8332 30072 8352
rect 29988 8324 30008 8332
rect 30016 8324 30044 8332
rect 30052 8324 30072 8332
rect 30108 8332 30192 8352
rect 30108 8324 30128 8332
rect 30136 8324 30164 8332
rect 30172 8324 30192 8332
rect 30228 8332 30312 8352
rect 30228 8324 30248 8332
rect 30256 8324 30284 8332
rect 30292 8324 30312 8332
rect 30348 8332 30432 8352
rect 30348 8324 30368 8332
rect 30376 8324 30404 8332
rect 30412 8324 30432 8332
rect 30468 8332 30552 8352
rect 30468 8324 30488 8332
rect 30496 8324 30524 8332
rect 30532 8324 30552 8332
rect 30588 8332 30672 8352
rect 30588 8324 30608 8332
rect 30616 8324 30644 8332
rect 30652 8324 30672 8332
rect 30708 8332 30792 8352
rect 30708 8324 30728 8332
rect 30736 8324 30764 8332
rect 30772 8324 30792 8332
rect 30828 8332 30912 8352
rect 30828 8324 30848 8332
rect 30856 8324 30884 8332
rect 30892 8324 30912 8332
rect 30948 8332 31032 8352
rect 30948 8324 30968 8332
rect 30976 8324 31004 8332
rect 31012 8324 31032 8332
rect 31068 8332 31152 8352
rect 31068 8324 31088 8332
rect 31096 8324 31124 8332
rect 31132 8324 31152 8332
rect 31188 8332 31272 8352
rect 31188 8324 31208 8332
rect 31216 8324 31244 8332
rect 31252 8324 31272 8332
rect 31308 8332 31392 8352
rect 31308 8324 31328 8332
rect 31336 8324 31364 8332
rect 31372 8324 31392 8332
rect 31428 8332 31512 8352
rect 31428 8324 31448 8332
rect 31456 8324 31484 8332
rect 31492 8324 31512 8332
rect 31548 8332 31632 8352
rect 31548 8324 31568 8332
rect 31576 8324 31604 8332
rect 31612 8324 31632 8332
rect 31668 8332 31752 8352
rect 31668 8324 31688 8332
rect 31696 8324 31724 8332
rect 31732 8324 31752 8332
rect 31788 8332 31872 8352
rect 31788 8324 31808 8332
rect 31816 8324 31844 8332
rect 31852 8324 31872 8332
rect 31908 8332 31992 8352
rect 31908 8324 31928 8332
rect 31936 8324 31964 8332
rect 31972 8324 31992 8332
rect 32028 8332 32112 8352
rect 32028 8324 32048 8332
rect 32056 8324 32084 8332
rect 32092 8324 32112 8332
rect 32148 8332 32232 8352
rect 32148 8324 32168 8332
rect 32176 8324 32204 8332
rect 32212 8324 32232 8332
rect 32268 8332 32352 8352
rect 32268 8324 32288 8332
rect 32296 8324 32324 8332
rect 32332 8324 32352 8332
rect 32388 8332 32472 8352
rect 32388 8324 32408 8332
rect 32416 8324 32444 8332
rect 32452 8324 32472 8332
rect 32508 8332 32592 8352
rect 32508 8324 32528 8332
rect 32536 8324 32564 8332
rect 32572 8324 32592 8332
rect 32628 8332 32712 8352
rect 32628 8324 32648 8332
rect 32656 8324 32684 8332
rect 32692 8324 32712 8332
rect 32748 8332 32832 8352
rect 32748 8324 32768 8332
rect 32776 8324 32804 8332
rect 32812 8324 32832 8332
rect 32868 8332 32952 8352
rect 32868 8324 32888 8332
rect 32896 8324 32924 8332
rect 32932 8324 32952 8332
rect 32988 8332 33072 8352
rect 32988 8324 33008 8332
rect 33016 8324 33044 8332
rect 33052 8324 33072 8332
rect 33108 8332 33192 8352
rect 33108 8324 33128 8332
rect 33136 8324 33164 8332
rect 33172 8324 33192 8332
rect 33228 8332 33312 8352
rect 33228 8324 33248 8332
rect 33256 8324 33284 8332
rect 33292 8324 33312 8332
rect 33348 8332 33432 8352
rect 33348 8324 33368 8332
rect 33376 8324 33404 8332
rect 33412 8324 33432 8332
rect 33468 8332 33552 8352
rect 33468 8324 33488 8332
rect 33496 8324 33524 8332
rect 33532 8324 33552 8332
rect 33588 8332 33672 8352
rect 33588 8324 33608 8332
rect 33616 8324 33644 8332
rect 33652 8324 33672 8332
rect 33708 8332 33792 8352
rect 33708 8324 33728 8332
rect 33736 8324 33764 8332
rect 33772 8324 33792 8332
rect 33828 8332 33912 8352
rect 33828 8324 33848 8332
rect 33856 8324 33884 8332
rect 33892 8324 33912 8332
rect 33948 8332 34032 8352
rect 33948 8324 33968 8332
rect 33976 8324 34004 8332
rect 34012 8324 34032 8332
rect 34068 8332 34152 8352
rect 34068 8324 34088 8332
rect 34096 8324 34124 8332
rect 34132 8324 34152 8332
rect 34188 8332 34272 8352
rect 34188 8324 34208 8332
rect 34216 8324 34244 8332
rect 34252 8324 34272 8332
rect 34308 8332 34392 8352
rect 34308 8324 34328 8332
rect 34336 8324 34364 8332
rect 34372 8324 34392 8332
rect 34428 8332 34512 8352
rect 34428 8324 34448 8332
rect 34456 8324 34484 8332
rect 34492 8324 34512 8332
rect 34548 8332 34632 8352
rect 34548 8324 34568 8332
rect 34576 8324 34604 8332
rect 34612 8324 34632 8332
rect 34668 8332 34752 8352
rect 34668 8324 34688 8332
rect 34696 8324 34724 8332
rect 34732 8324 34752 8332
rect 34788 8332 34872 8352
rect 34788 8324 34808 8332
rect 34816 8324 34844 8332
rect 34852 8324 34872 8332
rect 34908 8332 34992 8352
rect 34908 8324 34928 8332
rect 34936 8324 34964 8332
rect 34972 8324 34992 8332
rect 35028 8332 35112 8352
rect 35028 8324 35048 8332
rect 35056 8324 35084 8332
rect 35092 8324 35112 8332
rect 35148 8332 35232 8352
rect 35148 8324 35168 8332
rect 35176 8324 35204 8332
rect 35212 8324 35232 8332
rect 35268 8332 35352 8352
rect 35268 8324 35288 8332
rect 35296 8324 35324 8332
rect 35332 8324 35352 8332
rect 35388 8332 35472 8352
rect 35388 8324 35408 8332
rect 35416 8324 35444 8332
rect 35452 8324 35472 8332
rect 35508 8332 35592 8352
rect 35508 8324 35528 8332
rect 35536 8324 35564 8332
rect 35572 8324 35592 8332
rect 35628 8332 35712 8352
rect 35628 8324 35648 8332
rect 35656 8324 35684 8332
rect 35692 8324 35712 8332
rect 35748 8332 35832 8352
rect 35748 8324 35768 8332
rect 35776 8324 35804 8332
rect 35812 8324 35832 8332
rect 35868 8332 35952 8352
rect 35868 8324 35888 8332
rect 35896 8324 35924 8332
rect 35932 8324 35952 8332
rect 35988 8332 36072 8352
rect 35988 8324 36008 8332
rect 36016 8324 36044 8332
rect 36052 8324 36072 8332
rect 36108 8332 36192 8352
rect 36108 8324 36128 8332
rect 36136 8324 36164 8332
rect 36172 8324 36192 8332
rect 36228 8332 36312 8352
rect 36228 8324 36248 8332
rect 36256 8324 36284 8332
rect 36292 8324 36312 8332
rect 36348 8332 36432 8352
rect 36348 8324 36368 8332
rect 36376 8324 36404 8332
rect 36412 8324 36432 8332
rect 36468 8332 36552 8352
rect 36468 8324 36488 8332
rect 36496 8324 36524 8332
rect 36532 8324 36552 8332
rect 36588 8332 36672 8352
rect 36588 8324 36608 8332
rect 36616 8324 36644 8332
rect 36652 8324 36672 8332
rect 36708 8332 36792 8352
rect 36708 8324 36728 8332
rect 36736 8324 36764 8332
rect 36772 8324 36792 8332
rect 36828 8332 36912 8352
rect 36828 8324 36848 8332
rect 36856 8324 36884 8332
rect 36892 8324 36912 8332
rect 36948 8332 37032 8352
rect 36948 8324 36968 8332
rect 36976 8324 37004 8332
rect 37012 8324 37032 8332
rect 37068 8332 37152 8352
rect 37068 8324 37088 8332
rect 37096 8324 37124 8332
rect 37132 8324 37152 8332
rect 37188 8332 37272 8352
rect 37188 8324 37208 8332
rect 37216 8324 37244 8332
rect 37252 8324 37272 8332
rect 37308 8332 37392 8352
rect 37308 8324 37328 8332
rect 37336 8324 37364 8332
rect 37372 8324 37392 8332
rect 37428 8332 37512 8352
rect 37428 8324 37448 8332
rect 37456 8324 37484 8332
rect 37492 8324 37512 8332
rect 37548 8332 37632 8352
rect 37548 8324 37568 8332
rect 37576 8324 37604 8332
rect 37612 8324 37632 8332
rect 37668 8332 37752 8352
rect 37668 8324 37688 8332
rect 37696 8324 37724 8332
rect 37732 8324 37752 8332
rect 37788 8332 37872 8352
rect 37788 8324 37808 8332
rect 37816 8324 37844 8332
rect 37852 8324 37872 8332
rect 37908 8332 37992 8352
rect 37908 8324 37928 8332
rect 37936 8324 37964 8332
rect 37972 8324 37992 8332
rect 38028 8332 38112 8352
rect 38028 8324 38048 8332
rect 38056 8324 38084 8332
rect 38092 8324 38112 8332
rect 38148 8332 38232 8352
rect 38148 8324 38168 8332
rect 38176 8324 38204 8332
rect 38212 8324 38232 8332
rect 38268 8332 38352 8352
rect 38268 8324 38288 8332
rect 38296 8324 38324 8332
rect 38332 8324 38352 8332
rect 38388 8332 38472 8352
rect 38388 8324 38408 8332
rect 38416 8324 38444 8332
rect 38452 8324 38472 8332
rect 38508 8332 38592 8352
rect 38508 8324 38528 8332
rect 38536 8324 38564 8332
rect 38572 8324 38592 8332
rect 38628 8332 38712 8352
rect 38628 8324 38648 8332
rect 38656 8324 38684 8332
rect 38692 8324 38712 8332
rect 38748 8332 38832 8352
rect 38748 8324 38768 8332
rect 38776 8324 38804 8332
rect 38812 8324 38832 8332
rect 38868 8332 38952 8352
rect 38868 8324 38888 8332
rect 38896 8324 38924 8332
rect 38932 8324 38952 8332
rect 38988 8332 39072 8352
rect 38988 8324 39008 8332
rect 39016 8324 39044 8332
rect 39052 8324 39072 8332
rect 39108 8332 39192 8352
rect 39108 8324 39128 8332
rect 39136 8324 39164 8332
rect 39172 8324 39192 8332
rect 39228 8332 39312 8352
rect 39228 8324 39248 8332
rect 39256 8324 39284 8332
rect 39292 8324 39312 8332
rect 39348 8332 39432 8352
rect 39348 8324 39368 8332
rect 39376 8324 39404 8332
rect 39412 8324 39432 8332
rect 39468 8332 39552 8352
rect 39468 8324 39488 8332
rect 39496 8324 39524 8332
rect 39532 8324 39552 8332
rect 39588 8332 39672 8352
rect 39588 8324 39608 8332
rect 39616 8324 39644 8332
rect 39652 8324 39672 8332
rect 39708 8332 39792 8352
rect 39708 8324 39728 8332
rect 39736 8324 39764 8332
rect 39772 8324 39792 8332
rect 39828 8332 39912 8352
rect 39828 8324 39848 8332
rect 39856 8324 39884 8332
rect 39892 8324 39912 8332
rect 39948 8332 40032 8352
rect 39948 8324 39968 8332
rect 39976 8324 40004 8332
rect 40012 8324 40032 8332
rect 40068 8332 40152 8352
rect 40068 8324 40088 8332
rect 40096 8324 40124 8332
rect 40132 8324 40152 8332
rect 40188 8332 40272 8352
rect 40188 8324 40208 8332
rect 40216 8324 40244 8332
rect 40252 8324 40272 8332
rect 40308 8332 40392 8352
rect 40308 8324 40328 8332
rect 40336 8324 40364 8332
rect 40372 8324 40392 8332
rect 40428 8332 40512 8352
rect 40428 8324 40448 8332
rect 40456 8324 40484 8332
rect 40492 8324 40512 8332
rect 40548 8332 40632 8352
rect 40548 8324 40568 8332
rect 40576 8324 40604 8332
rect 40612 8324 40632 8332
rect 40668 8332 40752 8352
rect 40668 8324 40688 8332
rect 40696 8324 40724 8332
rect 40732 8324 40752 8332
rect 40788 8332 40872 8352
rect 40788 8324 40808 8332
rect 40816 8324 40844 8332
rect 40852 8324 40872 8332
rect 40908 8332 40992 8352
rect 40908 8324 40928 8332
rect 40936 8324 40964 8332
rect 40972 8324 40992 8332
rect 41028 8332 41112 8352
rect 41028 8324 41048 8332
rect 41056 8324 41084 8332
rect 41092 8324 41112 8332
rect 41148 8332 41232 8352
rect 41148 8324 41168 8332
rect 41176 8324 41204 8332
rect 41212 8324 41232 8332
rect 41268 8332 41352 8352
rect 41268 8324 41288 8332
rect 41296 8324 41324 8332
rect 41332 8324 41352 8332
rect 41388 8332 41472 8352
rect 41388 8324 41408 8332
rect 41416 8324 41444 8332
rect 41452 8324 41472 8332
rect 41508 8332 41592 8352
rect 41508 8324 41528 8332
rect 41536 8324 41564 8332
rect 41572 8324 41592 8332
rect 41628 8332 41712 8352
rect 41628 8324 41648 8332
rect 41656 8324 41684 8332
rect 41692 8324 41712 8332
rect 41748 8332 41832 8352
rect 41748 8324 41768 8332
rect 41776 8324 41804 8332
rect 41812 8324 41832 8332
rect 41868 8332 41952 8352
rect 41868 8324 41888 8332
rect 41896 8324 41924 8332
rect 41932 8324 41952 8332
rect 41988 8332 42072 8352
rect 41988 8324 42008 8332
rect 42016 8324 42044 8332
rect 42052 8324 42072 8332
rect 42108 8332 42192 8352
rect 42108 8324 42128 8332
rect 42136 8324 42164 8332
rect 42172 8324 42192 8332
rect 42228 8332 42312 8352
rect 42228 8324 42248 8332
rect 42256 8324 42284 8332
rect 42292 8324 42312 8332
rect 42348 8332 42432 8352
rect 42348 8324 42368 8332
rect 42376 8324 42404 8332
rect 42412 8324 42432 8332
rect 42468 8332 42552 8352
rect 42468 8324 42488 8332
rect 42496 8324 42524 8332
rect 42532 8324 42552 8332
rect 42588 8332 42672 8352
rect 42588 8324 42608 8332
rect 42616 8324 42644 8332
rect 42652 8324 42672 8332
rect 42708 8332 42792 8352
rect 42708 8324 42728 8332
rect 42736 8324 42764 8332
rect 42772 8324 42792 8332
rect 42828 8332 42912 8352
rect 42828 8324 42848 8332
rect 42856 8324 42884 8332
rect 42892 8324 42912 8332
rect 42948 8332 43032 8352
rect 42948 8324 42968 8332
rect 42976 8324 43004 8332
rect 43012 8324 43032 8332
rect 43068 8332 43152 8352
rect 43068 8324 43088 8332
rect 43096 8324 43124 8332
rect 43132 8324 43152 8332
rect 43188 8332 43272 8352
rect 43188 8324 43208 8332
rect 43216 8324 43244 8332
rect 43252 8324 43272 8332
rect 43308 8332 43392 8352
rect 43308 8324 43328 8332
rect 43336 8324 43364 8332
rect 43372 8324 43392 8332
rect 43428 8332 43512 8352
rect 43428 8324 43448 8332
rect 43456 8324 43484 8332
rect 43492 8324 43512 8332
rect 43548 8332 43632 8352
rect 43548 8324 43568 8332
rect 43576 8324 43604 8332
rect 43612 8324 43632 8332
rect 43668 8332 43752 8352
rect 43668 8324 43688 8332
rect 43696 8324 43724 8332
rect 43732 8324 43752 8332
rect 43788 8332 43872 8352
rect 43788 8324 43808 8332
rect 43816 8324 43844 8332
rect 43852 8324 43872 8332
rect 43908 8332 43992 8352
rect 43908 8324 43928 8332
rect 43936 8324 43964 8332
rect 43972 8324 43992 8332
rect 44028 8332 44112 8352
rect 44028 8324 44048 8332
rect 44056 8324 44084 8332
rect 44092 8324 44112 8332
rect 44148 8332 44232 8352
rect 44148 8324 44168 8332
rect 44176 8324 44204 8332
rect 44212 8324 44232 8332
rect 44268 8332 44352 8352
rect 44268 8324 44288 8332
rect 44296 8324 44324 8332
rect 44332 8324 44352 8332
rect 44388 8332 44472 8352
rect 44388 8324 44408 8332
rect 44416 8324 44444 8332
rect 44452 8324 44472 8332
rect 44508 8332 44592 8352
rect 44508 8324 44528 8332
rect 44536 8324 44564 8332
rect 44572 8324 44592 8332
rect 44628 8332 44712 8352
rect 44628 8324 44648 8332
rect 44656 8324 44684 8332
rect 44692 8324 44712 8332
rect 44748 8332 44832 8352
rect 44748 8324 44768 8332
rect 44776 8324 44804 8332
rect 44812 8324 44832 8332
rect 44868 8332 44952 8352
rect 44868 8324 44888 8332
rect 44896 8324 44924 8332
rect 44932 8324 44952 8332
rect 44988 8332 45072 8352
rect 44988 8324 45008 8332
rect 45016 8324 45044 8332
rect 45052 8324 45072 8332
rect 45108 8332 45192 8352
rect 45108 8324 45128 8332
rect 45136 8324 45164 8332
rect 45172 8324 45192 8332
rect 45228 8332 45312 8352
rect 45228 8324 45248 8332
rect 45256 8324 45284 8332
rect 45292 8324 45312 8332
rect 45348 8332 45432 8352
rect 45348 8324 45368 8332
rect 45376 8324 45404 8332
rect 45412 8324 45432 8332
rect 45468 8332 45552 8352
rect 45468 8324 45488 8332
rect 45496 8324 45524 8332
rect 45532 8324 45552 8332
rect 45588 8332 45672 8352
rect 45588 8324 45608 8332
rect 45616 8324 45644 8332
rect 45652 8324 45672 8332
rect 25936 8296 25992 8324
rect 26056 8296 26112 8324
rect 26176 8296 26232 8324
rect 26296 8296 26352 8324
rect 26416 8296 26472 8324
rect 26536 8296 26592 8324
rect 26656 8296 26712 8324
rect 26776 8296 26832 8324
rect 26896 8296 26952 8324
rect 27016 8296 27072 8324
rect 27136 8296 27192 8324
rect 27256 8296 27312 8324
rect 27376 8296 27432 8324
rect 27496 8296 27552 8324
rect 27616 8296 27672 8324
rect 27736 8296 27792 8324
rect 27856 8296 27912 8324
rect 27976 8296 28032 8324
rect 28096 8296 28152 8324
rect 28216 8296 28272 8324
rect 28336 8296 28392 8324
rect 28456 8296 28512 8324
rect 28576 8296 28632 8324
rect 28696 8296 28752 8324
rect 28816 8296 28872 8324
rect 28936 8296 28992 8324
rect 29056 8296 29112 8324
rect 29176 8296 29232 8324
rect 29296 8296 29352 8324
rect 29416 8296 29472 8324
rect 29536 8296 29592 8324
rect 29656 8296 29712 8324
rect 29776 8296 29832 8324
rect 29896 8296 29952 8324
rect 30016 8296 30072 8324
rect 30136 8296 30192 8324
rect 30256 8296 30312 8324
rect 30376 8296 30432 8324
rect 30496 8296 30552 8324
rect 30616 8296 30672 8324
rect 30736 8296 30792 8324
rect 30856 8296 30912 8324
rect 30976 8296 31032 8324
rect 31096 8296 31152 8324
rect 31216 8296 31272 8324
rect 31336 8296 31392 8324
rect 31456 8296 31512 8324
rect 31576 8296 31632 8324
rect 31696 8296 31752 8324
rect 31816 8296 31872 8324
rect 31936 8296 31992 8324
rect 32056 8296 32112 8324
rect 32176 8296 32232 8324
rect 32296 8296 32352 8324
rect 32416 8296 32472 8324
rect 32536 8296 32592 8324
rect 32656 8296 32712 8324
rect 32776 8296 32832 8324
rect 32896 8296 32952 8324
rect 33016 8296 33072 8324
rect 33136 8296 33192 8324
rect 33256 8296 33312 8324
rect 33376 8296 33432 8324
rect 33496 8296 33552 8324
rect 33616 8296 33672 8324
rect 33736 8296 33792 8324
rect 33856 8296 33912 8324
rect 33976 8296 34032 8324
rect 34096 8296 34152 8324
rect 34216 8296 34272 8324
rect 34336 8296 34392 8324
rect 34456 8296 34512 8324
rect 34576 8296 34632 8324
rect 34696 8296 34752 8324
rect 34816 8296 34872 8324
rect 34936 8296 34992 8324
rect 35056 8296 35112 8324
rect 35176 8296 35232 8324
rect 35296 8296 35352 8324
rect 35416 8296 35472 8324
rect 35536 8296 35592 8324
rect 35656 8296 35712 8324
rect 35776 8296 35832 8324
rect 35896 8296 35952 8324
rect 36016 8296 36072 8324
rect 36136 8296 36192 8324
rect 36256 8296 36312 8324
rect 36376 8296 36432 8324
rect 36496 8296 36552 8324
rect 36616 8296 36672 8324
rect 36736 8296 36792 8324
rect 36856 8296 36912 8324
rect 36976 8296 37032 8324
rect 37096 8296 37152 8324
rect 37216 8296 37272 8324
rect 37336 8296 37392 8324
rect 37456 8296 37512 8324
rect 37576 8296 37632 8324
rect 37696 8296 37752 8324
rect 37816 8296 37872 8324
rect 37936 8296 37992 8324
rect 38056 8296 38112 8324
rect 38176 8296 38232 8324
rect 38296 8296 38352 8324
rect 38416 8296 38472 8324
rect 38536 8296 38592 8324
rect 38656 8296 38712 8324
rect 38776 8296 38832 8324
rect 38896 8296 38952 8324
rect 39016 8296 39072 8324
rect 39136 8296 39192 8324
rect 39256 8296 39312 8324
rect 39376 8296 39432 8324
rect 39496 8296 39552 8324
rect 39616 8296 39672 8324
rect 39736 8296 39792 8324
rect 39856 8296 39912 8324
rect 39976 8296 40032 8324
rect 40096 8296 40152 8324
rect 40216 8296 40272 8324
rect 40336 8296 40392 8324
rect 40456 8296 40512 8324
rect 40576 8296 40632 8324
rect 40696 8296 40752 8324
rect 40816 8296 40872 8324
rect 40936 8296 40992 8324
rect 41056 8296 41112 8324
rect 41176 8296 41232 8324
rect 41296 8296 41352 8324
rect 41416 8296 41472 8324
rect 41536 8296 41592 8324
rect 41656 8296 41712 8324
rect 41776 8296 41832 8324
rect 41896 8296 41952 8324
rect 42016 8296 42072 8324
rect 42136 8296 42192 8324
rect 42256 8296 42312 8324
rect 42376 8296 42432 8324
rect 42496 8296 42552 8324
rect 42616 8296 42672 8324
rect 42736 8296 42792 8324
rect 42856 8296 42912 8324
rect 42976 8296 43032 8324
rect 43096 8296 43152 8324
rect 43216 8296 43272 8324
rect 43336 8296 43392 8324
rect 43456 8296 43512 8324
rect 43576 8296 43632 8324
rect 43696 8296 43752 8324
rect 43816 8296 43872 8324
rect 43936 8296 43992 8324
rect 44056 8296 44112 8324
rect 44176 8296 44232 8324
rect 44296 8296 44352 8324
rect 44416 8296 44472 8324
rect 44536 8296 44592 8324
rect 44656 8296 44712 8324
rect 44776 8296 44832 8324
rect 44896 8296 44952 8324
rect 45016 8296 45072 8324
rect 45136 8296 45192 8324
rect 45256 8296 45312 8324
rect 45376 8296 45432 8324
rect 45496 8296 45552 8324
rect 45616 8296 45672 8324
rect 25908 8152 25992 8172
rect 25908 8144 25928 8152
rect 25936 8144 25964 8152
rect 25972 8144 25992 8152
rect 26028 8152 26112 8172
rect 26028 8144 26048 8152
rect 26056 8144 26084 8152
rect 26092 8144 26112 8152
rect 26148 8152 26232 8172
rect 26148 8144 26168 8152
rect 26176 8144 26204 8152
rect 26212 8144 26232 8152
rect 26268 8152 26352 8172
rect 26268 8144 26288 8152
rect 26296 8144 26324 8152
rect 26332 8144 26352 8152
rect 26388 8152 26472 8172
rect 26388 8144 26408 8152
rect 26416 8144 26444 8152
rect 26452 8144 26472 8152
rect 26508 8152 26592 8172
rect 26508 8144 26528 8152
rect 26536 8144 26564 8152
rect 26572 8144 26592 8152
rect 26628 8152 26712 8172
rect 26628 8144 26648 8152
rect 26656 8144 26684 8152
rect 26692 8144 26712 8152
rect 26748 8152 26832 8172
rect 26748 8144 26768 8152
rect 26776 8144 26804 8152
rect 26812 8144 26832 8152
rect 26868 8152 26952 8172
rect 26868 8144 26888 8152
rect 26896 8144 26924 8152
rect 26932 8144 26952 8152
rect 26988 8152 27072 8172
rect 26988 8144 27008 8152
rect 27016 8144 27044 8152
rect 27052 8144 27072 8152
rect 27108 8152 27192 8172
rect 27108 8144 27128 8152
rect 27136 8144 27164 8152
rect 27172 8144 27192 8152
rect 27228 8152 27312 8172
rect 27228 8144 27248 8152
rect 27256 8144 27284 8152
rect 27292 8144 27312 8152
rect 27348 8152 27432 8172
rect 27348 8144 27368 8152
rect 27376 8144 27404 8152
rect 27412 8144 27432 8152
rect 27468 8152 27552 8172
rect 27468 8144 27488 8152
rect 27496 8144 27524 8152
rect 27532 8144 27552 8152
rect 27588 8152 27672 8172
rect 27588 8144 27608 8152
rect 27616 8144 27644 8152
rect 27652 8144 27672 8152
rect 27708 8152 27792 8172
rect 27708 8144 27728 8152
rect 27736 8144 27764 8152
rect 27772 8144 27792 8152
rect 27828 8152 27912 8172
rect 27828 8144 27848 8152
rect 27856 8144 27884 8152
rect 27892 8144 27912 8152
rect 27948 8152 28032 8172
rect 27948 8144 27968 8152
rect 27976 8144 28004 8152
rect 28012 8144 28032 8152
rect 28068 8152 28152 8172
rect 28068 8144 28088 8152
rect 28096 8144 28124 8152
rect 28132 8144 28152 8152
rect 28188 8152 28272 8172
rect 28188 8144 28208 8152
rect 28216 8144 28244 8152
rect 28252 8144 28272 8152
rect 28308 8152 28392 8172
rect 28308 8144 28328 8152
rect 28336 8144 28364 8152
rect 28372 8144 28392 8152
rect 28428 8152 28512 8172
rect 28428 8144 28448 8152
rect 28456 8144 28484 8152
rect 28492 8144 28512 8152
rect 28548 8152 28632 8172
rect 28548 8144 28568 8152
rect 28576 8144 28604 8152
rect 28612 8144 28632 8152
rect 28668 8152 28752 8172
rect 28668 8144 28688 8152
rect 28696 8144 28724 8152
rect 28732 8144 28752 8152
rect 28788 8152 28872 8172
rect 28788 8144 28808 8152
rect 28816 8144 28844 8152
rect 28852 8144 28872 8152
rect 28908 8152 28992 8172
rect 28908 8144 28928 8152
rect 28936 8144 28964 8152
rect 28972 8144 28992 8152
rect 29028 8152 29112 8172
rect 29028 8144 29048 8152
rect 29056 8144 29084 8152
rect 29092 8144 29112 8152
rect 29148 8152 29232 8172
rect 29148 8144 29168 8152
rect 29176 8144 29204 8152
rect 29212 8144 29232 8152
rect 29268 8152 29352 8172
rect 29268 8144 29288 8152
rect 29296 8144 29324 8152
rect 29332 8144 29352 8152
rect 29388 8152 29472 8172
rect 29388 8144 29408 8152
rect 29416 8144 29444 8152
rect 29452 8144 29472 8152
rect 29508 8152 29592 8172
rect 29508 8144 29528 8152
rect 29536 8144 29564 8152
rect 29572 8144 29592 8152
rect 29628 8152 29712 8172
rect 29628 8144 29648 8152
rect 29656 8144 29684 8152
rect 29692 8144 29712 8152
rect 29748 8152 29832 8172
rect 29748 8144 29768 8152
rect 29776 8144 29804 8152
rect 29812 8144 29832 8152
rect 29868 8152 29952 8172
rect 29868 8144 29888 8152
rect 29896 8144 29924 8152
rect 29932 8144 29952 8152
rect 29988 8152 30072 8172
rect 29988 8144 30008 8152
rect 30016 8144 30044 8152
rect 30052 8144 30072 8152
rect 30108 8152 30192 8172
rect 30108 8144 30128 8152
rect 30136 8144 30164 8152
rect 30172 8144 30192 8152
rect 30228 8152 30312 8172
rect 30228 8144 30248 8152
rect 30256 8144 30284 8152
rect 30292 8144 30312 8152
rect 30348 8152 30432 8172
rect 30348 8144 30368 8152
rect 30376 8144 30404 8152
rect 30412 8144 30432 8152
rect 30468 8152 30552 8172
rect 30468 8144 30488 8152
rect 30496 8144 30524 8152
rect 30532 8144 30552 8152
rect 30588 8152 30672 8172
rect 30588 8144 30608 8152
rect 30616 8144 30644 8152
rect 30652 8144 30672 8152
rect 30708 8152 30792 8172
rect 30708 8144 30728 8152
rect 30736 8144 30764 8152
rect 30772 8144 30792 8152
rect 30828 8152 30912 8172
rect 30828 8144 30848 8152
rect 30856 8144 30884 8152
rect 30892 8144 30912 8152
rect 30948 8152 31032 8172
rect 30948 8144 30968 8152
rect 30976 8144 31004 8152
rect 31012 8144 31032 8152
rect 31068 8152 31152 8172
rect 31068 8144 31088 8152
rect 31096 8144 31124 8152
rect 31132 8144 31152 8152
rect 31188 8152 31272 8172
rect 31188 8144 31208 8152
rect 31216 8144 31244 8152
rect 31252 8144 31272 8152
rect 31308 8152 31392 8172
rect 31308 8144 31328 8152
rect 31336 8144 31364 8152
rect 31372 8144 31392 8152
rect 31428 8152 31512 8172
rect 31428 8144 31448 8152
rect 31456 8144 31484 8152
rect 31492 8144 31512 8152
rect 31548 8152 31632 8172
rect 31548 8144 31568 8152
rect 31576 8144 31604 8152
rect 31612 8144 31632 8152
rect 31668 8152 31752 8172
rect 31668 8144 31688 8152
rect 31696 8144 31724 8152
rect 31732 8144 31752 8152
rect 31788 8152 31872 8172
rect 31788 8144 31808 8152
rect 31816 8144 31844 8152
rect 31852 8144 31872 8152
rect 31908 8152 31992 8172
rect 31908 8144 31928 8152
rect 31936 8144 31964 8152
rect 31972 8144 31992 8152
rect 32028 8152 32112 8172
rect 32028 8144 32048 8152
rect 32056 8144 32084 8152
rect 32092 8144 32112 8152
rect 32148 8152 32232 8172
rect 32148 8144 32168 8152
rect 32176 8144 32204 8152
rect 32212 8144 32232 8152
rect 32268 8152 32352 8172
rect 32268 8144 32288 8152
rect 32296 8144 32324 8152
rect 32332 8144 32352 8152
rect 32388 8152 32472 8172
rect 32388 8144 32408 8152
rect 32416 8144 32444 8152
rect 32452 8144 32472 8152
rect 32508 8152 32592 8172
rect 32508 8144 32528 8152
rect 32536 8144 32564 8152
rect 32572 8144 32592 8152
rect 32628 8152 32712 8172
rect 32628 8144 32648 8152
rect 32656 8144 32684 8152
rect 32692 8144 32712 8152
rect 32748 8152 32832 8172
rect 32748 8144 32768 8152
rect 32776 8144 32804 8152
rect 32812 8144 32832 8152
rect 32868 8152 32952 8172
rect 32868 8144 32888 8152
rect 32896 8144 32924 8152
rect 32932 8144 32952 8152
rect 32988 8152 33072 8172
rect 32988 8144 33008 8152
rect 33016 8144 33044 8152
rect 33052 8144 33072 8152
rect 33108 8152 33192 8172
rect 33108 8144 33128 8152
rect 33136 8144 33164 8152
rect 33172 8144 33192 8152
rect 33228 8152 33312 8172
rect 33228 8144 33248 8152
rect 33256 8144 33284 8152
rect 33292 8144 33312 8152
rect 33348 8152 33432 8172
rect 33348 8144 33368 8152
rect 33376 8144 33404 8152
rect 33412 8144 33432 8152
rect 33468 8152 33552 8172
rect 33468 8144 33488 8152
rect 33496 8144 33524 8152
rect 33532 8144 33552 8152
rect 33588 8152 33672 8172
rect 33588 8144 33608 8152
rect 33616 8144 33644 8152
rect 33652 8144 33672 8152
rect 33708 8152 33792 8172
rect 33708 8144 33728 8152
rect 33736 8144 33764 8152
rect 33772 8144 33792 8152
rect 33828 8152 33912 8172
rect 33828 8144 33848 8152
rect 33856 8144 33884 8152
rect 33892 8144 33912 8152
rect 33948 8152 34032 8172
rect 33948 8144 33968 8152
rect 33976 8144 34004 8152
rect 34012 8144 34032 8152
rect 34068 8152 34152 8172
rect 34068 8144 34088 8152
rect 34096 8144 34124 8152
rect 34132 8144 34152 8152
rect 34188 8152 34272 8172
rect 34188 8144 34208 8152
rect 34216 8144 34244 8152
rect 34252 8144 34272 8152
rect 34308 8152 34392 8172
rect 34308 8144 34328 8152
rect 34336 8144 34364 8152
rect 34372 8144 34392 8152
rect 34428 8152 34512 8172
rect 34428 8144 34448 8152
rect 34456 8144 34484 8152
rect 34492 8144 34512 8152
rect 34548 8152 34632 8172
rect 34548 8144 34568 8152
rect 34576 8144 34604 8152
rect 34612 8144 34632 8152
rect 34668 8152 34752 8172
rect 34668 8144 34688 8152
rect 34696 8144 34724 8152
rect 34732 8144 34752 8152
rect 34788 8152 34872 8172
rect 34788 8144 34808 8152
rect 34816 8144 34844 8152
rect 34852 8144 34872 8152
rect 34908 8152 34992 8172
rect 34908 8144 34928 8152
rect 34936 8144 34964 8152
rect 34972 8144 34992 8152
rect 35028 8152 35112 8172
rect 35028 8144 35048 8152
rect 35056 8144 35084 8152
rect 35092 8144 35112 8152
rect 35148 8152 35232 8172
rect 35148 8144 35168 8152
rect 35176 8144 35204 8152
rect 35212 8144 35232 8152
rect 35268 8152 35352 8172
rect 35268 8144 35288 8152
rect 35296 8144 35324 8152
rect 35332 8144 35352 8152
rect 35388 8152 35472 8172
rect 35388 8144 35408 8152
rect 35416 8144 35444 8152
rect 35452 8144 35472 8152
rect 35508 8152 35592 8172
rect 35508 8144 35528 8152
rect 35536 8144 35564 8152
rect 35572 8144 35592 8152
rect 35628 8152 35712 8172
rect 35628 8144 35648 8152
rect 35656 8144 35684 8152
rect 35692 8144 35712 8152
rect 35748 8152 35832 8172
rect 35748 8144 35768 8152
rect 35776 8144 35804 8152
rect 35812 8144 35832 8152
rect 35868 8152 35952 8172
rect 35868 8144 35888 8152
rect 35896 8144 35924 8152
rect 35932 8144 35952 8152
rect 35988 8152 36072 8172
rect 35988 8144 36008 8152
rect 36016 8144 36044 8152
rect 36052 8144 36072 8152
rect 36108 8152 36192 8172
rect 36108 8144 36128 8152
rect 36136 8144 36164 8152
rect 36172 8144 36192 8152
rect 36228 8152 36312 8172
rect 36228 8144 36248 8152
rect 36256 8144 36284 8152
rect 36292 8144 36312 8152
rect 36348 8152 36432 8172
rect 36348 8144 36368 8152
rect 36376 8144 36404 8152
rect 36412 8144 36432 8152
rect 36468 8152 36552 8172
rect 36468 8144 36488 8152
rect 36496 8144 36524 8152
rect 36532 8144 36552 8152
rect 36588 8152 36672 8172
rect 36588 8144 36608 8152
rect 36616 8144 36644 8152
rect 36652 8144 36672 8152
rect 36708 8152 36792 8172
rect 36708 8144 36728 8152
rect 36736 8144 36764 8152
rect 36772 8144 36792 8152
rect 36828 8152 36912 8172
rect 36828 8144 36848 8152
rect 36856 8144 36884 8152
rect 36892 8144 36912 8152
rect 36948 8152 37032 8172
rect 36948 8144 36968 8152
rect 36976 8144 37004 8152
rect 37012 8144 37032 8152
rect 37068 8152 37152 8172
rect 37068 8144 37088 8152
rect 37096 8144 37124 8152
rect 37132 8144 37152 8152
rect 37188 8152 37272 8172
rect 37188 8144 37208 8152
rect 37216 8144 37244 8152
rect 37252 8144 37272 8152
rect 37308 8152 37392 8172
rect 37308 8144 37328 8152
rect 37336 8144 37364 8152
rect 37372 8144 37392 8152
rect 37428 8152 37512 8172
rect 37428 8144 37448 8152
rect 37456 8144 37484 8152
rect 37492 8144 37512 8152
rect 37548 8152 37632 8172
rect 37548 8144 37568 8152
rect 37576 8144 37604 8152
rect 37612 8144 37632 8152
rect 37668 8152 37752 8172
rect 37668 8144 37688 8152
rect 37696 8144 37724 8152
rect 37732 8144 37752 8152
rect 37788 8152 37872 8172
rect 37788 8144 37808 8152
rect 37816 8144 37844 8152
rect 37852 8144 37872 8152
rect 37908 8152 37992 8172
rect 37908 8144 37928 8152
rect 37936 8144 37964 8152
rect 37972 8144 37992 8152
rect 38028 8152 38112 8172
rect 38028 8144 38048 8152
rect 38056 8144 38084 8152
rect 38092 8144 38112 8152
rect 38148 8152 38232 8172
rect 38148 8144 38168 8152
rect 38176 8144 38204 8152
rect 38212 8144 38232 8152
rect 38268 8152 38352 8172
rect 38268 8144 38288 8152
rect 38296 8144 38324 8152
rect 38332 8144 38352 8152
rect 38388 8152 38472 8172
rect 38388 8144 38408 8152
rect 38416 8144 38444 8152
rect 38452 8144 38472 8152
rect 38508 8152 38592 8172
rect 38508 8144 38528 8152
rect 38536 8144 38564 8152
rect 38572 8144 38592 8152
rect 38628 8152 38712 8172
rect 38628 8144 38648 8152
rect 38656 8144 38684 8152
rect 38692 8144 38712 8152
rect 38748 8152 38832 8172
rect 38748 8144 38768 8152
rect 38776 8144 38804 8152
rect 38812 8144 38832 8152
rect 38868 8152 38952 8172
rect 38868 8144 38888 8152
rect 38896 8144 38924 8152
rect 38932 8144 38952 8152
rect 38988 8152 39072 8172
rect 38988 8144 39008 8152
rect 39016 8144 39044 8152
rect 39052 8144 39072 8152
rect 39108 8152 39192 8172
rect 39108 8144 39128 8152
rect 39136 8144 39164 8152
rect 39172 8144 39192 8152
rect 39228 8152 39312 8172
rect 39228 8144 39248 8152
rect 39256 8144 39284 8152
rect 39292 8144 39312 8152
rect 39348 8152 39432 8172
rect 39348 8144 39368 8152
rect 39376 8144 39404 8152
rect 39412 8144 39432 8152
rect 39468 8152 39552 8172
rect 39468 8144 39488 8152
rect 39496 8144 39524 8152
rect 39532 8144 39552 8152
rect 39588 8152 39672 8172
rect 39588 8144 39608 8152
rect 39616 8144 39644 8152
rect 39652 8144 39672 8152
rect 39708 8152 39792 8172
rect 39708 8144 39728 8152
rect 39736 8144 39764 8152
rect 39772 8144 39792 8152
rect 39828 8152 39912 8172
rect 39828 8144 39848 8152
rect 39856 8144 39884 8152
rect 39892 8144 39912 8152
rect 39948 8152 40032 8172
rect 39948 8144 39968 8152
rect 39976 8144 40004 8152
rect 40012 8144 40032 8152
rect 40068 8152 40152 8172
rect 40068 8144 40088 8152
rect 40096 8144 40124 8152
rect 40132 8144 40152 8152
rect 40188 8152 40272 8172
rect 40188 8144 40208 8152
rect 40216 8144 40244 8152
rect 40252 8144 40272 8152
rect 40308 8152 40392 8172
rect 40308 8144 40328 8152
rect 40336 8144 40364 8152
rect 40372 8144 40392 8152
rect 40428 8152 40512 8172
rect 40428 8144 40448 8152
rect 40456 8144 40484 8152
rect 40492 8144 40512 8152
rect 40548 8152 40632 8172
rect 40548 8144 40568 8152
rect 40576 8144 40604 8152
rect 40612 8144 40632 8152
rect 40668 8152 40752 8172
rect 40668 8144 40688 8152
rect 40696 8144 40724 8152
rect 40732 8144 40752 8152
rect 40788 8152 40872 8172
rect 40788 8144 40808 8152
rect 40816 8144 40844 8152
rect 40852 8144 40872 8152
rect 40908 8152 40992 8172
rect 40908 8144 40928 8152
rect 40936 8144 40964 8152
rect 40972 8144 40992 8152
rect 41028 8152 41112 8172
rect 41028 8144 41048 8152
rect 41056 8144 41084 8152
rect 41092 8144 41112 8152
rect 41148 8152 41232 8172
rect 41148 8144 41168 8152
rect 41176 8144 41204 8152
rect 41212 8144 41232 8152
rect 41268 8152 41352 8172
rect 41268 8144 41288 8152
rect 41296 8144 41324 8152
rect 41332 8144 41352 8152
rect 41388 8152 41472 8172
rect 41388 8144 41408 8152
rect 41416 8144 41444 8152
rect 41452 8144 41472 8152
rect 41508 8152 41592 8172
rect 41508 8144 41528 8152
rect 41536 8144 41564 8152
rect 41572 8144 41592 8152
rect 41628 8152 41712 8172
rect 41628 8144 41648 8152
rect 41656 8144 41684 8152
rect 41692 8144 41712 8152
rect 41748 8152 41832 8172
rect 41748 8144 41768 8152
rect 41776 8144 41804 8152
rect 41812 8144 41832 8152
rect 41868 8152 41952 8172
rect 41868 8144 41888 8152
rect 41896 8144 41924 8152
rect 41932 8144 41952 8152
rect 41988 8152 42072 8172
rect 41988 8144 42008 8152
rect 42016 8144 42044 8152
rect 42052 8144 42072 8152
rect 42108 8152 42192 8172
rect 42108 8144 42128 8152
rect 42136 8144 42164 8152
rect 42172 8144 42192 8152
rect 42228 8152 42312 8172
rect 42228 8144 42248 8152
rect 42256 8144 42284 8152
rect 42292 8144 42312 8152
rect 42348 8152 42432 8172
rect 42348 8144 42368 8152
rect 42376 8144 42404 8152
rect 42412 8144 42432 8152
rect 42468 8152 42552 8172
rect 42468 8144 42488 8152
rect 42496 8144 42524 8152
rect 42532 8144 42552 8152
rect 42588 8152 42672 8172
rect 42588 8144 42608 8152
rect 42616 8144 42644 8152
rect 42652 8144 42672 8152
rect 42708 8152 42792 8172
rect 42708 8144 42728 8152
rect 42736 8144 42764 8152
rect 42772 8144 42792 8152
rect 42828 8152 42912 8172
rect 42828 8144 42848 8152
rect 42856 8144 42884 8152
rect 42892 8144 42912 8152
rect 42948 8152 43032 8172
rect 42948 8144 42968 8152
rect 42976 8144 43004 8152
rect 43012 8144 43032 8152
rect 43068 8152 43152 8172
rect 43068 8144 43088 8152
rect 43096 8144 43124 8152
rect 43132 8144 43152 8152
rect 43188 8152 43272 8172
rect 43188 8144 43208 8152
rect 43216 8144 43244 8152
rect 43252 8144 43272 8152
rect 43308 8152 43392 8172
rect 43308 8144 43328 8152
rect 43336 8144 43364 8152
rect 43372 8144 43392 8152
rect 43428 8152 43512 8172
rect 43428 8144 43448 8152
rect 43456 8144 43484 8152
rect 43492 8144 43512 8152
rect 43548 8152 43632 8172
rect 43548 8144 43568 8152
rect 43576 8144 43604 8152
rect 43612 8144 43632 8152
rect 43668 8152 43752 8172
rect 43668 8144 43688 8152
rect 43696 8144 43724 8152
rect 43732 8144 43752 8152
rect 43788 8152 43872 8172
rect 43788 8144 43808 8152
rect 43816 8144 43844 8152
rect 43852 8144 43872 8152
rect 43908 8152 43992 8172
rect 43908 8144 43928 8152
rect 43936 8144 43964 8152
rect 43972 8144 43992 8152
rect 44028 8152 44112 8172
rect 44028 8144 44048 8152
rect 44056 8144 44084 8152
rect 44092 8144 44112 8152
rect 44148 8152 44232 8172
rect 44148 8144 44168 8152
rect 44176 8144 44204 8152
rect 44212 8144 44232 8152
rect 44268 8152 44352 8172
rect 44268 8144 44288 8152
rect 44296 8144 44324 8152
rect 44332 8144 44352 8152
rect 44388 8152 44472 8172
rect 44388 8144 44408 8152
rect 44416 8144 44444 8152
rect 44452 8144 44472 8152
rect 44508 8152 44592 8172
rect 44508 8144 44528 8152
rect 44536 8144 44564 8152
rect 44572 8144 44592 8152
rect 44628 8152 44712 8172
rect 44628 8144 44648 8152
rect 44656 8144 44684 8152
rect 44692 8144 44712 8152
rect 44748 8152 44832 8172
rect 44748 8144 44768 8152
rect 44776 8144 44804 8152
rect 44812 8144 44832 8152
rect 44868 8152 44952 8172
rect 44868 8144 44888 8152
rect 44896 8144 44924 8152
rect 44932 8144 44952 8152
rect 44988 8152 45072 8172
rect 44988 8144 45008 8152
rect 45016 8144 45044 8152
rect 45052 8144 45072 8152
rect 45108 8152 45192 8172
rect 45108 8144 45128 8152
rect 45136 8144 45164 8152
rect 45172 8144 45192 8152
rect 45228 8152 45312 8172
rect 45228 8144 45248 8152
rect 45256 8144 45284 8152
rect 45292 8144 45312 8152
rect 45348 8152 45432 8172
rect 45348 8144 45368 8152
rect 45376 8144 45404 8152
rect 45412 8144 45432 8152
rect 45468 8152 45552 8172
rect 45468 8144 45488 8152
rect 45496 8144 45524 8152
rect 45532 8144 45552 8152
rect 45588 8152 45672 8172
rect 45588 8144 45608 8152
rect 45616 8144 45644 8152
rect 45652 8144 45672 8152
rect 25936 8116 25992 8144
rect 26056 8116 26112 8144
rect 26176 8116 26232 8144
rect 26296 8116 26352 8144
rect 26416 8116 26472 8144
rect 26536 8116 26592 8144
rect 26656 8116 26712 8144
rect 26776 8116 26832 8144
rect 26896 8116 26952 8144
rect 27016 8116 27072 8144
rect 27136 8116 27192 8144
rect 27256 8116 27312 8144
rect 27376 8116 27432 8144
rect 27496 8116 27552 8144
rect 27616 8116 27672 8144
rect 27736 8116 27792 8144
rect 27856 8116 27912 8144
rect 27976 8116 28032 8144
rect 28096 8116 28152 8144
rect 28216 8116 28272 8144
rect 28336 8116 28392 8144
rect 28456 8116 28512 8144
rect 28576 8116 28632 8144
rect 28696 8116 28752 8144
rect 28816 8116 28872 8144
rect 28936 8116 28992 8144
rect 29056 8116 29112 8144
rect 29176 8116 29232 8144
rect 29296 8116 29352 8144
rect 29416 8116 29472 8144
rect 29536 8116 29592 8144
rect 29656 8116 29712 8144
rect 29776 8116 29832 8144
rect 29896 8116 29952 8144
rect 30016 8116 30072 8144
rect 30136 8116 30192 8144
rect 30256 8116 30312 8144
rect 30376 8116 30432 8144
rect 30496 8116 30552 8144
rect 30616 8116 30672 8144
rect 30736 8116 30792 8144
rect 30856 8116 30912 8144
rect 30976 8116 31032 8144
rect 31096 8116 31152 8144
rect 31216 8116 31272 8144
rect 31336 8116 31392 8144
rect 31456 8116 31512 8144
rect 31576 8116 31632 8144
rect 31696 8116 31752 8144
rect 31816 8116 31872 8144
rect 31936 8116 31992 8144
rect 32056 8116 32112 8144
rect 32176 8116 32232 8144
rect 32296 8116 32352 8144
rect 32416 8116 32472 8144
rect 32536 8116 32592 8144
rect 32656 8116 32712 8144
rect 32776 8116 32832 8144
rect 32896 8116 32952 8144
rect 33016 8116 33072 8144
rect 33136 8116 33192 8144
rect 33256 8116 33312 8144
rect 33376 8116 33432 8144
rect 33496 8116 33552 8144
rect 33616 8116 33672 8144
rect 33736 8116 33792 8144
rect 33856 8116 33912 8144
rect 33976 8116 34032 8144
rect 34096 8116 34152 8144
rect 34216 8116 34272 8144
rect 34336 8116 34392 8144
rect 34456 8116 34512 8144
rect 34576 8116 34632 8144
rect 34696 8116 34752 8144
rect 34816 8116 34872 8144
rect 34936 8116 34992 8144
rect 35056 8116 35112 8144
rect 35176 8116 35232 8144
rect 35296 8116 35352 8144
rect 35416 8116 35472 8144
rect 35536 8116 35592 8144
rect 35656 8116 35712 8144
rect 35776 8116 35832 8144
rect 35896 8116 35952 8144
rect 36016 8116 36072 8144
rect 36136 8116 36192 8144
rect 36256 8116 36312 8144
rect 36376 8116 36432 8144
rect 36496 8116 36552 8144
rect 36616 8116 36672 8144
rect 36736 8116 36792 8144
rect 36856 8116 36912 8144
rect 36976 8116 37032 8144
rect 37096 8116 37152 8144
rect 37216 8116 37272 8144
rect 37336 8116 37392 8144
rect 37456 8116 37512 8144
rect 37576 8116 37632 8144
rect 37696 8116 37752 8144
rect 37816 8116 37872 8144
rect 37936 8116 37992 8144
rect 38056 8116 38112 8144
rect 38176 8116 38232 8144
rect 38296 8116 38352 8144
rect 38416 8116 38472 8144
rect 38536 8116 38592 8144
rect 38656 8116 38712 8144
rect 38776 8116 38832 8144
rect 38896 8116 38952 8144
rect 39016 8116 39072 8144
rect 39136 8116 39192 8144
rect 39256 8116 39312 8144
rect 39376 8116 39432 8144
rect 39496 8116 39552 8144
rect 39616 8116 39672 8144
rect 39736 8116 39792 8144
rect 39856 8116 39912 8144
rect 39976 8116 40032 8144
rect 40096 8116 40152 8144
rect 40216 8116 40272 8144
rect 40336 8116 40392 8144
rect 40456 8116 40512 8144
rect 40576 8116 40632 8144
rect 40696 8116 40752 8144
rect 40816 8116 40872 8144
rect 40936 8116 40992 8144
rect 41056 8116 41112 8144
rect 41176 8116 41232 8144
rect 41296 8116 41352 8144
rect 41416 8116 41472 8144
rect 41536 8116 41592 8144
rect 41656 8116 41712 8144
rect 41776 8116 41832 8144
rect 41896 8116 41952 8144
rect 42016 8116 42072 8144
rect 42136 8116 42192 8144
rect 42256 8116 42312 8144
rect 42376 8116 42432 8144
rect 42496 8116 42552 8144
rect 42616 8116 42672 8144
rect 42736 8116 42792 8144
rect 42856 8116 42912 8144
rect 42976 8116 43032 8144
rect 43096 8116 43152 8144
rect 43216 8116 43272 8144
rect 43336 8116 43392 8144
rect 43456 8116 43512 8144
rect 43576 8116 43632 8144
rect 43696 8116 43752 8144
rect 43816 8116 43872 8144
rect 43936 8116 43992 8144
rect 44056 8116 44112 8144
rect 44176 8116 44232 8144
rect 44296 8116 44352 8144
rect 44416 8116 44472 8144
rect 44536 8116 44592 8144
rect 44656 8116 44712 8144
rect 44776 8116 44832 8144
rect 44896 8116 44952 8144
rect 45016 8116 45072 8144
rect 45136 8116 45192 8144
rect 45256 8116 45312 8144
rect 45376 8116 45432 8144
rect 45496 8116 45552 8144
rect 45616 8116 45672 8144
rect 25908 7972 25992 7992
rect 25908 7964 25928 7972
rect 25936 7964 25964 7972
rect 25972 7964 25992 7972
rect 26028 7972 26112 7992
rect 26028 7964 26048 7972
rect 26056 7964 26084 7972
rect 26092 7964 26112 7972
rect 26148 7972 26232 7992
rect 26148 7964 26168 7972
rect 26176 7964 26204 7972
rect 26212 7964 26232 7972
rect 26268 7972 26352 7992
rect 26268 7964 26288 7972
rect 26296 7964 26324 7972
rect 26332 7964 26352 7972
rect 26388 7972 26472 7992
rect 26388 7964 26408 7972
rect 26416 7964 26444 7972
rect 26452 7964 26472 7972
rect 26508 7972 26592 7992
rect 26508 7964 26528 7972
rect 26536 7964 26564 7972
rect 26572 7964 26592 7972
rect 26628 7972 26712 7992
rect 26628 7964 26648 7972
rect 26656 7964 26684 7972
rect 26692 7964 26712 7972
rect 26748 7972 26832 7992
rect 26748 7964 26768 7972
rect 26776 7964 26804 7972
rect 26812 7964 26832 7972
rect 26868 7972 26952 7992
rect 26868 7964 26888 7972
rect 26896 7964 26924 7972
rect 26932 7964 26952 7972
rect 26988 7972 27072 7992
rect 26988 7964 27008 7972
rect 27016 7964 27044 7972
rect 27052 7964 27072 7972
rect 27108 7972 27192 7992
rect 27108 7964 27128 7972
rect 27136 7964 27164 7972
rect 27172 7964 27192 7972
rect 27228 7972 27312 7992
rect 27228 7964 27248 7972
rect 27256 7964 27284 7972
rect 27292 7964 27312 7972
rect 27348 7972 27432 7992
rect 27348 7964 27368 7972
rect 27376 7964 27404 7972
rect 27412 7964 27432 7972
rect 27468 7972 27552 7992
rect 27468 7964 27488 7972
rect 27496 7964 27524 7972
rect 27532 7964 27552 7972
rect 27588 7972 27672 7992
rect 27588 7964 27608 7972
rect 27616 7964 27644 7972
rect 27652 7964 27672 7972
rect 27708 7972 27792 7992
rect 27708 7964 27728 7972
rect 27736 7964 27764 7972
rect 27772 7964 27792 7972
rect 27828 7972 27912 7992
rect 27828 7964 27848 7972
rect 27856 7964 27884 7972
rect 27892 7964 27912 7972
rect 27948 7972 28032 7992
rect 27948 7964 27968 7972
rect 27976 7964 28004 7972
rect 28012 7964 28032 7972
rect 28068 7972 28152 7992
rect 28068 7964 28088 7972
rect 28096 7964 28124 7972
rect 28132 7964 28152 7972
rect 28188 7972 28272 7992
rect 28188 7964 28208 7972
rect 28216 7964 28244 7972
rect 28252 7964 28272 7972
rect 28308 7972 28392 7992
rect 28308 7964 28328 7972
rect 28336 7964 28364 7972
rect 28372 7964 28392 7972
rect 28428 7972 28512 7992
rect 28428 7964 28448 7972
rect 28456 7964 28484 7972
rect 28492 7964 28512 7972
rect 28548 7972 28632 7992
rect 28548 7964 28568 7972
rect 28576 7964 28604 7972
rect 28612 7964 28632 7972
rect 28668 7972 28752 7992
rect 28668 7964 28688 7972
rect 28696 7964 28724 7972
rect 28732 7964 28752 7972
rect 28788 7972 28872 7992
rect 28788 7964 28808 7972
rect 28816 7964 28844 7972
rect 28852 7964 28872 7972
rect 28908 7972 28992 7992
rect 28908 7964 28928 7972
rect 28936 7964 28964 7972
rect 28972 7964 28992 7972
rect 29028 7972 29112 7992
rect 29028 7964 29048 7972
rect 29056 7964 29084 7972
rect 29092 7964 29112 7972
rect 29148 7972 29232 7992
rect 29148 7964 29168 7972
rect 29176 7964 29204 7972
rect 29212 7964 29232 7972
rect 29268 7972 29352 7992
rect 29268 7964 29288 7972
rect 29296 7964 29324 7972
rect 29332 7964 29352 7972
rect 29388 7972 29472 7992
rect 29388 7964 29408 7972
rect 29416 7964 29444 7972
rect 29452 7964 29472 7972
rect 29508 7972 29592 7992
rect 29508 7964 29528 7972
rect 29536 7964 29564 7972
rect 29572 7964 29592 7972
rect 29628 7972 29712 7992
rect 29628 7964 29648 7972
rect 29656 7964 29684 7972
rect 29692 7964 29712 7972
rect 29748 7972 29832 7992
rect 29748 7964 29768 7972
rect 29776 7964 29804 7972
rect 29812 7964 29832 7972
rect 29868 7972 29952 7992
rect 29868 7964 29888 7972
rect 29896 7964 29924 7972
rect 29932 7964 29952 7972
rect 29988 7972 30072 7992
rect 29988 7964 30008 7972
rect 30016 7964 30044 7972
rect 30052 7964 30072 7972
rect 30108 7972 30192 7992
rect 30108 7964 30128 7972
rect 30136 7964 30164 7972
rect 30172 7964 30192 7972
rect 30228 7972 30312 7992
rect 30228 7964 30248 7972
rect 30256 7964 30284 7972
rect 30292 7964 30312 7972
rect 30348 7972 30432 7992
rect 30348 7964 30368 7972
rect 30376 7964 30404 7972
rect 30412 7964 30432 7972
rect 30468 7972 30552 7992
rect 30468 7964 30488 7972
rect 30496 7964 30524 7972
rect 30532 7964 30552 7972
rect 30588 7972 30672 7992
rect 30588 7964 30608 7972
rect 30616 7964 30644 7972
rect 30652 7964 30672 7972
rect 30708 7972 30792 7992
rect 30708 7964 30728 7972
rect 30736 7964 30764 7972
rect 30772 7964 30792 7972
rect 30828 7972 30912 7992
rect 30828 7964 30848 7972
rect 30856 7964 30884 7972
rect 30892 7964 30912 7972
rect 30948 7972 31032 7992
rect 30948 7964 30968 7972
rect 30976 7964 31004 7972
rect 31012 7964 31032 7972
rect 31068 7972 31152 7992
rect 31068 7964 31088 7972
rect 31096 7964 31124 7972
rect 31132 7964 31152 7972
rect 31188 7972 31272 7992
rect 31188 7964 31208 7972
rect 31216 7964 31244 7972
rect 31252 7964 31272 7972
rect 31308 7972 31392 7992
rect 31308 7964 31328 7972
rect 31336 7964 31364 7972
rect 31372 7964 31392 7972
rect 31428 7972 31512 7992
rect 31428 7964 31448 7972
rect 31456 7964 31484 7972
rect 31492 7964 31512 7972
rect 31548 7972 31632 7992
rect 31548 7964 31568 7972
rect 31576 7964 31604 7972
rect 31612 7964 31632 7972
rect 31668 7972 31752 7992
rect 31668 7964 31688 7972
rect 31696 7964 31724 7972
rect 31732 7964 31752 7972
rect 31788 7972 31872 7992
rect 31788 7964 31808 7972
rect 31816 7964 31844 7972
rect 31852 7964 31872 7972
rect 31908 7972 31992 7992
rect 31908 7964 31928 7972
rect 31936 7964 31964 7972
rect 31972 7964 31992 7972
rect 32028 7972 32112 7992
rect 32028 7964 32048 7972
rect 32056 7964 32084 7972
rect 32092 7964 32112 7972
rect 32148 7972 32232 7992
rect 32148 7964 32168 7972
rect 32176 7964 32204 7972
rect 32212 7964 32232 7972
rect 32268 7972 32352 7992
rect 32268 7964 32288 7972
rect 32296 7964 32324 7972
rect 32332 7964 32352 7972
rect 32388 7972 32472 7992
rect 32388 7964 32408 7972
rect 32416 7964 32444 7972
rect 32452 7964 32472 7972
rect 32508 7972 32592 7992
rect 32508 7964 32528 7972
rect 32536 7964 32564 7972
rect 32572 7964 32592 7972
rect 32628 7972 32712 7992
rect 32628 7964 32648 7972
rect 32656 7964 32684 7972
rect 32692 7964 32712 7972
rect 32748 7972 32832 7992
rect 32748 7964 32768 7972
rect 32776 7964 32804 7972
rect 32812 7964 32832 7972
rect 32868 7972 32952 7992
rect 32868 7964 32888 7972
rect 32896 7964 32924 7972
rect 32932 7964 32952 7972
rect 32988 7972 33072 7992
rect 32988 7964 33008 7972
rect 33016 7964 33044 7972
rect 33052 7964 33072 7972
rect 33108 7972 33192 7992
rect 33108 7964 33128 7972
rect 33136 7964 33164 7972
rect 33172 7964 33192 7972
rect 33228 7972 33312 7992
rect 33228 7964 33248 7972
rect 33256 7964 33284 7972
rect 33292 7964 33312 7972
rect 33348 7972 33432 7992
rect 33348 7964 33368 7972
rect 33376 7964 33404 7972
rect 33412 7964 33432 7972
rect 33468 7972 33552 7992
rect 33468 7964 33488 7972
rect 33496 7964 33524 7972
rect 33532 7964 33552 7972
rect 33588 7972 33672 7992
rect 33588 7964 33608 7972
rect 33616 7964 33644 7972
rect 33652 7964 33672 7972
rect 33708 7972 33792 7992
rect 33708 7964 33728 7972
rect 33736 7964 33764 7972
rect 33772 7964 33792 7972
rect 33828 7972 33912 7992
rect 33828 7964 33848 7972
rect 33856 7964 33884 7972
rect 33892 7964 33912 7972
rect 33948 7972 34032 7992
rect 33948 7964 33968 7972
rect 33976 7964 34004 7972
rect 34012 7964 34032 7972
rect 34068 7972 34152 7992
rect 34068 7964 34088 7972
rect 34096 7964 34124 7972
rect 34132 7964 34152 7972
rect 34188 7972 34272 7992
rect 34188 7964 34208 7972
rect 34216 7964 34244 7972
rect 34252 7964 34272 7972
rect 34308 7972 34392 7992
rect 34308 7964 34328 7972
rect 34336 7964 34364 7972
rect 34372 7964 34392 7972
rect 34428 7972 34512 7992
rect 34428 7964 34448 7972
rect 34456 7964 34484 7972
rect 34492 7964 34512 7972
rect 34548 7972 34632 7992
rect 34548 7964 34568 7972
rect 34576 7964 34604 7972
rect 34612 7964 34632 7972
rect 34668 7972 34752 7992
rect 34668 7964 34688 7972
rect 34696 7964 34724 7972
rect 34732 7964 34752 7972
rect 34788 7972 34872 7992
rect 34788 7964 34808 7972
rect 34816 7964 34844 7972
rect 34852 7964 34872 7972
rect 34908 7972 34992 7992
rect 34908 7964 34928 7972
rect 34936 7964 34964 7972
rect 34972 7964 34992 7972
rect 35028 7972 35112 7992
rect 35028 7964 35048 7972
rect 35056 7964 35084 7972
rect 35092 7964 35112 7972
rect 35148 7972 35232 7992
rect 35148 7964 35168 7972
rect 35176 7964 35204 7972
rect 35212 7964 35232 7972
rect 35268 7972 35352 7992
rect 35268 7964 35288 7972
rect 35296 7964 35324 7972
rect 35332 7964 35352 7972
rect 35388 7972 35472 7992
rect 35388 7964 35408 7972
rect 35416 7964 35444 7972
rect 35452 7964 35472 7972
rect 35508 7972 35592 7992
rect 35508 7964 35528 7972
rect 35536 7964 35564 7972
rect 35572 7964 35592 7972
rect 35628 7972 35712 7992
rect 35628 7964 35648 7972
rect 35656 7964 35684 7972
rect 35692 7964 35712 7972
rect 35748 7972 35832 7992
rect 35748 7964 35768 7972
rect 35776 7964 35804 7972
rect 35812 7964 35832 7972
rect 35868 7972 35952 7992
rect 35868 7964 35888 7972
rect 35896 7964 35924 7972
rect 35932 7964 35952 7972
rect 35988 7972 36072 7992
rect 35988 7964 36008 7972
rect 36016 7964 36044 7972
rect 36052 7964 36072 7972
rect 36108 7972 36192 7992
rect 36108 7964 36128 7972
rect 36136 7964 36164 7972
rect 36172 7964 36192 7972
rect 36228 7972 36312 7992
rect 36228 7964 36248 7972
rect 36256 7964 36284 7972
rect 36292 7964 36312 7972
rect 36348 7972 36432 7992
rect 36348 7964 36368 7972
rect 36376 7964 36404 7972
rect 36412 7964 36432 7972
rect 36468 7972 36552 7992
rect 36468 7964 36488 7972
rect 36496 7964 36524 7972
rect 36532 7964 36552 7972
rect 36588 7972 36672 7992
rect 36588 7964 36608 7972
rect 36616 7964 36644 7972
rect 36652 7964 36672 7972
rect 36708 7972 36792 7992
rect 36708 7964 36728 7972
rect 36736 7964 36764 7972
rect 36772 7964 36792 7972
rect 36828 7972 36912 7992
rect 36828 7964 36848 7972
rect 36856 7964 36884 7972
rect 36892 7964 36912 7972
rect 36948 7972 37032 7992
rect 36948 7964 36968 7972
rect 36976 7964 37004 7972
rect 37012 7964 37032 7972
rect 37068 7972 37152 7992
rect 37068 7964 37088 7972
rect 37096 7964 37124 7972
rect 37132 7964 37152 7972
rect 37188 7972 37272 7992
rect 37188 7964 37208 7972
rect 37216 7964 37244 7972
rect 37252 7964 37272 7972
rect 37308 7972 37392 7992
rect 37308 7964 37328 7972
rect 37336 7964 37364 7972
rect 37372 7964 37392 7972
rect 37428 7972 37512 7992
rect 37428 7964 37448 7972
rect 37456 7964 37484 7972
rect 37492 7964 37512 7972
rect 37548 7972 37632 7992
rect 37548 7964 37568 7972
rect 37576 7964 37604 7972
rect 37612 7964 37632 7972
rect 37668 7972 37752 7992
rect 37668 7964 37688 7972
rect 37696 7964 37724 7972
rect 37732 7964 37752 7972
rect 37788 7972 37872 7992
rect 37788 7964 37808 7972
rect 37816 7964 37844 7972
rect 37852 7964 37872 7972
rect 37908 7972 37992 7992
rect 37908 7964 37928 7972
rect 37936 7964 37964 7972
rect 37972 7964 37992 7972
rect 38028 7972 38112 7992
rect 38028 7964 38048 7972
rect 38056 7964 38084 7972
rect 38092 7964 38112 7972
rect 38148 7972 38232 7992
rect 38148 7964 38168 7972
rect 38176 7964 38204 7972
rect 38212 7964 38232 7972
rect 38268 7972 38352 7992
rect 38268 7964 38288 7972
rect 38296 7964 38324 7972
rect 38332 7964 38352 7972
rect 38388 7972 38472 7992
rect 38388 7964 38408 7972
rect 38416 7964 38444 7972
rect 38452 7964 38472 7972
rect 38508 7972 38592 7992
rect 38508 7964 38528 7972
rect 38536 7964 38564 7972
rect 38572 7964 38592 7972
rect 38628 7972 38712 7992
rect 38628 7964 38648 7972
rect 38656 7964 38684 7972
rect 38692 7964 38712 7972
rect 38748 7972 38832 7992
rect 38748 7964 38768 7972
rect 38776 7964 38804 7972
rect 38812 7964 38832 7972
rect 38868 7972 38952 7992
rect 38868 7964 38888 7972
rect 38896 7964 38924 7972
rect 38932 7964 38952 7972
rect 38988 7972 39072 7992
rect 38988 7964 39008 7972
rect 39016 7964 39044 7972
rect 39052 7964 39072 7972
rect 39108 7972 39192 7992
rect 39108 7964 39128 7972
rect 39136 7964 39164 7972
rect 39172 7964 39192 7972
rect 39228 7972 39312 7992
rect 39228 7964 39248 7972
rect 39256 7964 39284 7972
rect 39292 7964 39312 7972
rect 39348 7972 39432 7992
rect 39348 7964 39368 7972
rect 39376 7964 39404 7972
rect 39412 7964 39432 7972
rect 39468 7972 39552 7992
rect 39468 7964 39488 7972
rect 39496 7964 39524 7972
rect 39532 7964 39552 7972
rect 39588 7972 39672 7992
rect 39588 7964 39608 7972
rect 39616 7964 39644 7972
rect 39652 7964 39672 7972
rect 39708 7972 39792 7992
rect 39708 7964 39728 7972
rect 39736 7964 39764 7972
rect 39772 7964 39792 7972
rect 39828 7972 39912 7992
rect 39828 7964 39848 7972
rect 39856 7964 39884 7972
rect 39892 7964 39912 7972
rect 39948 7972 40032 7992
rect 39948 7964 39968 7972
rect 39976 7964 40004 7972
rect 40012 7964 40032 7972
rect 40068 7972 40152 7992
rect 40068 7964 40088 7972
rect 40096 7964 40124 7972
rect 40132 7964 40152 7972
rect 40188 7972 40272 7992
rect 40188 7964 40208 7972
rect 40216 7964 40244 7972
rect 40252 7964 40272 7972
rect 40308 7972 40392 7992
rect 40308 7964 40328 7972
rect 40336 7964 40364 7972
rect 40372 7964 40392 7972
rect 40428 7972 40512 7992
rect 40428 7964 40448 7972
rect 40456 7964 40484 7972
rect 40492 7964 40512 7972
rect 40548 7972 40632 7992
rect 40548 7964 40568 7972
rect 40576 7964 40604 7972
rect 40612 7964 40632 7972
rect 40668 7972 40752 7992
rect 40668 7964 40688 7972
rect 40696 7964 40724 7972
rect 40732 7964 40752 7972
rect 40788 7972 40872 7992
rect 40788 7964 40808 7972
rect 40816 7964 40844 7972
rect 40852 7964 40872 7972
rect 40908 7972 40992 7992
rect 40908 7964 40928 7972
rect 40936 7964 40964 7972
rect 40972 7964 40992 7972
rect 41028 7972 41112 7992
rect 41028 7964 41048 7972
rect 41056 7964 41084 7972
rect 41092 7964 41112 7972
rect 41148 7972 41232 7992
rect 41148 7964 41168 7972
rect 41176 7964 41204 7972
rect 41212 7964 41232 7972
rect 41268 7972 41352 7992
rect 41268 7964 41288 7972
rect 41296 7964 41324 7972
rect 41332 7964 41352 7972
rect 41388 7972 41472 7992
rect 41388 7964 41408 7972
rect 41416 7964 41444 7972
rect 41452 7964 41472 7972
rect 41508 7972 41592 7992
rect 41508 7964 41528 7972
rect 41536 7964 41564 7972
rect 41572 7964 41592 7972
rect 41628 7972 41712 7992
rect 41628 7964 41648 7972
rect 41656 7964 41684 7972
rect 41692 7964 41712 7972
rect 41748 7972 41832 7992
rect 41748 7964 41768 7972
rect 41776 7964 41804 7972
rect 41812 7964 41832 7972
rect 41868 7972 41952 7992
rect 41868 7964 41888 7972
rect 41896 7964 41924 7972
rect 41932 7964 41952 7972
rect 41988 7972 42072 7992
rect 41988 7964 42008 7972
rect 42016 7964 42044 7972
rect 42052 7964 42072 7972
rect 42108 7972 42192 7992
rect 42108 7964 42128 7972
rect 42136 7964 42164 7972
rect 42172 7964 42192 7972
rect 42228 7972 42312 7992
rect 42228 7964 42248 7972
rect 42256 7964 42284 7972
rect 42292 7964 42312 7972
rect 42348 7972 42432 7992
rect 42348 7964 42368 7972
rect 42376 7964 42404 7972
rect 42412 7964 42432 7972
rect 42468 7972 42552 7992
rect 42468 7964 42488 7972
rect 42496 7964 42524 7972
rect 42532 7964 42552 7972
rect 42588 7972 42672 7992
rect 42588 7964 42608 7972
rect 42616 7964 42644 7972
rect 42652 7964 42672 7972
rect 42708 7972 42792 7992
rect 42708 7964 42728 7972
rect 42736 7964 42764 7972
rect 42772 7964 42792 7972
rect 42828 7972 42912 7992
rect 42828 7964 42848 7972
rect 42856 7964 42884 7972
rect 42892 7964 42912 7972
rect 42948 7972 43032 7992
rect 42948 7964 42968 7972
rect 42976 7964 43004 7972
rect 43012 7964 43032 7972
rect 43068 7972 43152 7992
rect 43068 7964 43088 7972
rect 43096 7964 43124 7972
rect 43132 7964 43152 7972
rect 43188 7972 43272 7992
rect 43188 7964 43208 7972
rect 43216 7964 43244 7972
rect 43252 7964 43272 7972
rect 43308 7972 43392 7992
rect 43308 7964 43328 7972
rect 43336 7964 43364 7972
rect 43372 7964 43392 7972
rect 43428 7972 43512 7992
rect 43428 7964 43448 7972
rect 43456 7964 43484 7972
rect 43492 7964 43512 7972
rect 43548 7972 43632 7992
rect 43548 7964 43568 7972
rect 43576 7964 43604 7972
rect 43612 7964 43632 7972
rect 43668 7972 43752 7992
rect 43668 7964 43688 7972
rect 43696 7964 43724 7972
rect 43732 7964 43752 7972
rect 43788 7972 43872 7992
rect 43788 7964 43808 7972
rect 43816 7964 43844 7972
rect 43852 7964 43872 7972
rect 43908 7972 43992 7992
rect 43908 7964 43928 7972
rect 43936 7964 43964 7972
rect 43972 7964 43992 7972
rect 44028 7972 44112 7992
rect 44028 7964 44048 7972
rect 44056 7964 44084 7972
rect 44092 7964 44112 7972
rect 44148 7972 44232 7992
rect 44148 7964 44168 7972
rect 44176 7964 44204 7972
rect 44212 7964 44232 7972
rect 44268 7972 44352 7992
rect 44268 7964 44288 7972
rect 44296 7964 44324 7972
rect 44332 7964 44352 7972
rect 44388 7972 44472 7992
rect 44388 7964 44408 7972
rect 44416 7964 44444 7972
rect 44452 7964 44472 7972
rect 44508 7972 44592 7992
rect 44508 7964 44528 7972
rect 44536 7964 44564 7972
rect 44572 7964 44592 7972
rect 44628 7972 44712 7992
rect 44628 7964 44648 7972
rect 44656 7964 44684 7972
rect 44692 7964 44712 7972
rect 44748 7972 44832 7992
rect 44748 7964 44768 7972
rect 44776 7964 44804 7972
rect 44812 7964 44832 7972
rect 44868 7972 44952 7992
rect 44868 7964 44888 7972
rect 44896 7964 44924 7972
rect 44932 7964 44952 7972
rect 44988 7972 45072 7992
rect 44988 7964 45008 7972
rect 45016 7964 45044 7972
rect 45052 7964 45072 7972
rect 45108 7972 45192 7992
rect 45108 7964 45128 7972
rect 45136 7964 45164 7972
rect 45172 7964 45192 7972
rect 45228 7972 45312 7992
rect 45228 7964 45248 7972
rect 45256 7964 45284 7972
rect 45292 7964 45312 7972
rect 45348 7972 45432 7992
rect 45348 7964 45368 7972
rect 45376 7964 45404 7972
rect 45412 7964 45432 7972
rect 45468 7972 45552 7992
rect 45468 7964 45488 7972
rect 45496 7964 45524 7972
rect 45532 7964 45552 7972
rect 45588 7972 45672 7992
rect 45588 7964 45608 7972
rect 45616 7964 45644 7972
rect 45652 7964 45672 7972
rect 25936 7936 25992 7964
rect 26056 7936 26112 7964
rect 26176 7936 26232 7964
rect 26296 7936 26352 7964
rect 26416 7936 26472 7964
rect 26536 7936 26592 7964
rect 26656 7936 26712 7964
rect 26776 7936 26832 7964
rect 26896 7936 26952 7964
rect 27016 7936 27072 7964
rect 27136 7936 27192 7964
rect 27256 7936 27312 7964
rect 27376 7936 27432 7964
rect 27496 7936 27552 7964
rect 27616 7936 27672 7964
rect 27736 7936 27792 7964
rect 27856 7936 27912 7964
rect 27976 7936 28032 7964
rect 28096 7936 28152 7964
rect 28216 7936 28272 7964
rect 28336 7936 28392 7964
rect 28456 7936 28512 7964
rect 28576 7936 28632 7964
rect 28696 7936 28752 7964
rect 28816 7936 28872 7964
rect 28936 7936 28992 7964
rect 29056 7936 29112 7964
rect 29176 7936 29232 7964
rect 29296 7936 29352 7964
rect 29416 7936 29472 7964
rect 29536 7936 29592 7964
rect 29656 7936 29712 7964
rect 29776 7936 29832 7964
rect 29896 7936 29952 7964
rect 30016 7936 30072 7964
rect 30136 7936 30192 7964
rect 30256 7936 30312 7964
rect 30376 7936 30432 7964
rect 30496 7936 30552 7964
rect 30616 7936 30672 7964
rect 30736 7936 30792 7964
rect 30856 7936 30912 7964
rect 30976 7936 31032 7964
rect 31096 7936 31152 7964
rect 31216 7936 31272 7964
rect 31336 7936 31392 7964
rect 31456 7936 31512 7964
rect 31576 7936 31632 7964
rect 31696 7936 31752 7964
rect 31816 7936 31872 7964
rect 31936 7936 31992 7964
rect 32056 7936 32112 7964
rect 32176 7936 32232 7964
rect 32296 7936 32352 7964
rect 32416 7936 32472 7964
rect 32536 7936 32592 7964
rect 32656 7936 32712 7964
rect 32776 7936 32832 7964
rect 32896 7936 32952 7964
rect 33016 7936 33072 7964
rect 33136 7936 33192 7964
rect 33256 7936 33312 7964
rect 33376 7936 33432 7964
rect 33496 7936 33552 7964
rect 33616 7936 33672 7964
rect 33736 7936 33792 7964
rect 33856 7936 33912 7964
rect 33976 7936 34032 7964
rect 34096 7936 34152 7964
rect 34216 7936 34272 7964
rect 34336 7936 34392 7964
rect 34456 7936 34512 7964
rect 34576 7936 34632 7964
rect 34696 7936 34752 7964
rect 34816 7936 34872 7964
rect 34936 7936 34992 7964
rect 35056 7936 35112 7964
rect 35176 7936 35232 7964
rect 35296 7936 35352 7964
rect 35416 7936 35472 7964
rect 35536 7936 35592 7964
rect 35656 7936 35712 7964
rect 35776 7936 35832 7964
rect 35896 7936 35952 7964
rect 36016 7936 36072 7964
rect 36136 7936 36192 7964
rect 36256 7936 36312 7964
rect 36376 7936 36432 7964
rect 36496 7936 36552 7964
rect 36616 7936 36672 7964
rect 36736 7936 36792 7964
rect 36856 7936 36912 7964
rect 36976 7936 37032 7964
rect 37096 7936 37152 7964
rect 37216 7936 37272 7964
rect 37336 7936 37392 7964
rect 37456 7936 37512 7964
rect 37576 7936 37632 7964
rect 37696 7936 37752 7964
rect 37816 7936 37872 7964
rect 37936 7936 37992 7964
rect 38056 7936 38112 7964
rect 38176 7936 38232 7964
rect 38296 7936 38352 7964
rect 38416 7936 38472 7964
rect 38536 7936 38592 7964
rect 38656 7936 38712 7964
rect 38776 7936 38832 7964
rect 38896 7936 38952 7964
rect 39016 7936 39072 7964
rect 39136 7936 39192 7964
rect 39256 7936 39312 7964
rect 39376 7936 39432 7964
rect 39496 7936 39552 7964
rect 39616 7936 39672 7964
rect 39736 7936 39792 7964
rect 39856 7936 39912 7964
rect 39976 7936 40032 7964
rect 40096 7936 40152 7964
rect 40216 7936 40272 7964
rect 40336 7936 40392 7964
rect 40456 7936 40512 7964
rect 40576 7936 40632 7964
rect 40696 7936 40752 7964
rect 40816 7936 40872 7964
rect 40936 7936 40992 7964
rect 41056 7936 41112 7964
rect 41176 7936 41232 7964
rect 41296 7936 41352 7964
rect 41416 7936 41472 7964
rect 41536 7936 41592 7964
rect 41656 7936 41712 7964
rect 41776 7936 41832 7964
rect 41896 7936 41952 7964
rect 42016 7936 42072 7964
rect 42136 7936 42192 7964
rect 42256 7936 42312 7964
rect 42376 7936 42432 7964
rect 42496 7936 42552 7964
rect 42616 7936 42672 7964
rect 42736 7936 42792 7964
rect 42856 7936 42912 7964
rect 42976 7936 43032 7964
rect 43096 7936 43152 7964
rect 43216 7936 43272 7964
rect 43336 7936 43392 7964
rect 43456 7936 43512 7964
rect 43576 7936 43632 7964
rect 43696 7936 43752 7964
rect 43816 7936 43872 7964
rect 43936 7936 43992 7964
rect 44056 7936 44112 7964
rect 44176 7936 44232 7964
rect 44296 7936 44352 7964
rect 44416 7936 44472 7964
rect 44536 7936 44592 7964
rect 44656 7936 44712 7964
rect 44776 7936 44832 7964
rect 44896 7936 44952 7964
rect 45016 7936 45072 7964
rect 45136 7936 45192 7964
rect 45256 7936 45312 7964
rect 45376 7936 45432 7964
rect 45496 7936 45552 7964
rect 45616 7936 45672 7964
rect 25908 7792 25992 7812
rect 25908 7784 25928 7792
rect 25936 7784 25964 7792
rect 25972 7784 25992 7792
rect 26028 7792 26112 7812
rect 26028 7784 26048 7792
rect 26056 7784 26084 7792
rect 26092 7784 26112 7792
rect 26148 7792 26232 7812
rect 26148 7784 26168 7792
rect 26176 7784 26204 7792
rect 26212 7784 26232 7792
rect 26268 7792 26352 7812
rect 26268 7784 26288 7792
rect 26296 7784 26324 7792
rect 26332 7784 26352 7792
rect 26388 7792 26472 7812
rect 26388 7784 26408 7792
rect 26416 7784 26444 7792
rect 26452 7784 26472 7792
rect 26508 7792 26592 7812
rect 26508 7784 26528 7792
rect 26536 7784 26564 7792
rect 26572 7784 26592 7792
rect 26628 7792 26712 7812
rect 26628 7784 26648 7792
rect 26656 7784 26684 7792
rect 26692 7784 26712 7792
rect 26748 7792 26832 7812
rect 26748 7784 26768 7792
rect 26776 7784 26804 7792
rect 26812 7784 26832 7792
rect 26868 7792 26952 7812
rect 26868 7784 26888 7792
rect 26896 7784 26924 7792
rect 26932 7784 26952 7792
rect 26988 7792 27072 7812
rect 26988 7784 27008 7792
rect 27016 7784 27044 7792
rect 27052 7784 27072 7792
rect 27108 7792 27192 7812
rect 27108 7784 27128 7792
rect 27136 7784 27164 7792
rect 27172 7784 27192 7792
rect 27228 7792 27312 7812
rect 27228 7784 27248 7792
rect 27256 7784 27284 7792
rect 27292 7784 27312 7792
rect 27348 7792 27432 7812
rect 27348 7784 27368 7792
rect 27376 7784 27404 7792
rect 27412 7784 27432 7792
rect 27468 7792 27552 7812
rect 27468 7784 27488 7792
rect 27496 7784 27524 7792
rect 27532 7784 27552 7792
rect 27588 7792 27672 7812
rect 27588 7784 27608 7792
rect 27616 7784 27644 7792
rect 27652 7784 27672 7792
rect 27708 7792 27792 7812
rect 27708 7784 27728 7792
rect 27736 7784 27764 7792
rect 27772 7784 27792 7792
rect 27828 7792 27912 7812
rect 27828 7784 27848 7792
rect 27856 7784 27884 7792
rect 27892 7784 27912 7792
rect 27948 7792 28032 7812
rect 27948 7784 27968 7792
rect 27976 7784 28004 7792
rect 28012 7784 28032 7792
rect 28068 7792 28152 7812
rect 28068 7784 28088 7792
rect 28096 7784 28124 7792
rect 28132 7784 28152 7792
rect 28188 7792 28272 7812
rect 28188 7784 28208 7792
rect 28216 7784 28244 7792
rect 28252 7784 28272 7792
rect 28308 7792 28392 7812
rect 28308 7784 28328 7792
rect 28336 7784 28364 7792
rect 28372 7784 28392 7792
rect 28428 7792 28512 7812
rect 28428 7784 28448 7792
rect 28456 7784 28484 7792
rect 28492 7784 28512 7792
rect 28548 7792 28632 7812
rect 28548 7784 28568 7792
rect 28576 7784 28604 7792
rect 28612 7784 28632 7792
rect 28668 7792 28752 7812
rect 28668 7784 28688 7792
rect 28696 7784 28724 7792
rect 28732 7784 28752 7792
rect 28788 7792 28872 7812
rect 28788 7784 28808 7792
rect 28816 7784 28844 7792
rect 28852 7784 28872 7792
rect 28908 7792 28992 7812
rect 28908 7784 28928 7792
rect 28936 7784 28964 7792
rect 28972 7784 28992 7792
rect 29028 7792 29112 7812
rect 29028 7784 29048 7792
rect 29056 7784 29084 7792
rect 29092 7784 29112 7792
rect 29148 7792 29232 7812
rect 29148 7784 29168 7792
rect 29176 7784 29204 7792
rect 29212 7784 29232 7792
rect 29268 7792 29352 7812
rect 29268 7784 29288 7792
rect 29296 7784 29324 7792
rect 29332 7784 29352 7792
rect 29388 7792 29472 7812
rect 29388 7784 29408 7792
rect 29416 7784 29444 7792
rect 29452 7784 29472 7792
rect 29508 7792 29592 7812
rect 29508 7784 29528 7792
rect 29536 7784 29564 7792
rect 29572 7784 29592 7792
rect 29628 7792 29712 7812
rect 29628 7784 29648 7792
rect 29656 7784 29684 7792
rect 29692 7784 29712 7792
rect 29748 7792 29832 7812
rect 29748 7784 29768 7792
rect 29776 7784 29804 7792
rect 29812 7784 29832 7792
rect 29868 7792 29952 7812
rect 29868 7784 29888 7792
rect 29896 7784 29924 7792
rect 29932 7784 29952 7792
rect 29988 7792 30072 7812
rect 29988 7784 30008 7792
rect 30016 7784 30044 7792
rect 30052 7784 30072 7792
rect 30108 7792 30192 7812
rect 30108 7784 30128 7792
rect 30136 7784 30164 7792
rect 30172 7784 30192 7792
rect 30228 7792 30312 7812
rect 30228 7784 30248 7792
rect 30256 7784 30284 7792
rect 30292 7784 30312 7792
rect 30348 7792 30432 7812
rect 30348 7784 30368 7792
rect 30376 7784 30404 7792
rect 30412 7784 30432 7792
rect 30468 7792 30552 7812
rect 30468 7784 30488 7792
rect 30496 7784 30524 7792
rect 30532 7784 30552 7792
rect 30588 7792 30672 7812
rect 30588 7784 30608 7792
rect 30616 7784 30644 7792
rect 30652 7784 30672 7792
rect 30708 7792 30792 7812
rect 30708 7784 30728 7792
rect 30736 7784 30764 7792
rect 30772 7784 30792 7792
rect 30828 7792 30912 7812
rect 30828 7784 30848 7792
rect 30856 7784 30884 7792
rect 30892 7784 30912 7792
rect 30948 7792 31032 7812
rect 30948 7784 30968 7792
rect 30976 7784 31004 7792
rect 31012 7784 31032 7792
rect 31068 7792 31152 7812
rect 31068 7784 31088 7792
rect 31096 7784 31124 7792
rect 31132 7784 31152 7792
rect 31188 7792 31272 7812
rect 31188 7784 31208 7792
rect 31216 7784 31244 7792
rect 31252 7784 31272 7792
rect 31308 7792 31392 7812
rect 31308 7784 31328 7792
rect 31336 7784 31364 7792
rect 31372 7784 31392 7792
rect 31428 7792 31512 7812
rect 31428 7784 31448 7792
rect 31456 7784 31484 7792
rect 31492 7784 31512 7792
rect 31548 7792 31632 7812
rect 31548 7784 31568 7792
rect 31576 7784 31604 7792
rect 31612 7784 31632 7792
rect 31668 7792 31752 7812
rect 31668 7784 31688 7792
rect 31696 7784 31724 7792
rect 31732 7784 31752 7792
rect 31788 7792 31872 7812
rect 31788 7784 31808 7792
rect 31816 7784 31844 7792
rect 31852 7784 31872 7792
rect 31908 7792 31992 7812
rect 31908 7784 31928 7792
rect 31936 7784 31964 7792
rect 31972 7784 31992 7792
rect 32028 7792 32112 7812
rect 32028 7784 32048 7792
rect 32056 7784 32084 7792
rect 32092 7784 32112 7792
rect 32148 7792 32232 7812
rect 32148 7784 32168 7792
rect 32176 7784 32204 7792
rect 32212 7784 32232 7792
rect 32268 7792 32352 7812
rect 32268 7784 32288 7792
rect 32296 7784 32324 7792
rect 32332 7784 32352 7792
rect 32388 7792 32472 7812
rect 32388 7784 32408 7792
rect 32416 7784 32444 7792
rect 32452 7784 32472 7792
rect 32508 7792 32592 7812
rect 32508 7784 32528 7792
rect 32536 7784 32564 7792
rect 32572 7784 32592 7792
rect 32628 7792 32712 7812
rect 32628 7784 32648 7792
rect 32656 7784 32684 7792
rect 32692 7784 32712 7792
rect 32748 7792 32832 7812
rect 32748 7784 32768 7792
rect 32776 7784 32804 7792
rect 32812 7784 32832 7792
rect 32868 7792 32952 7812
rect 32868 7784 32888 7792
rect 32896 7784 32924 7792
rect 32932 7784 32952 7792
rect 32988 7792 33072 7812
rect 32988 7784 33008 7792
rect 33016 7784 33044 7792
rect 33052 7784 33072 7792
rect 33108 7792 33192 7812
rect 33108 7784 33128 7792
rect 33136 7784 33164 7792
rect 33172 7784 33192 7792
rect 33228 7792 33312 7812
rect 33228 7784 33248 7792
rect 33256 7784 33284 7792
rect 33292 7784 33312 7792
rect 33348 7792 33432 7812
rect 33348 7784 33368 7792
rect 33376 7784 33404 7792
rect 33412 7784 33432 7792
rect 33468 7792 33552 7812
rect 33468 7784 33488 7792
rect 33496 7784 33524 7792
rect 33532 7784 33552 7792
rect 33588 7792 33672 7812
rect 33588 7784 33608 7792
rect 33616 7784 33644 7792
rect 33652 7784 33672 7792
rect 33708 7792 33792 7812
rect 33708 7784 33728 7792
rect 33736 7784 33764 7792
rect 33772 7784 33792 7792
rect 33828 7792 33912 7812
rect 33828 7784 33848 7792
rect 33856 7784 33884 7792
rect 33892 7784 33912 7792
rect 33948 7792 34032 7812
rect 33948 7784 33968 7792
rect 33976 7784 34004 7792
rect 34012 7784 34032 7792
rect 34068 7792 34152 7812
rect 34068 7784 34088 7792
rect 34096 7784 34124 7792
rect 34132 7784 34152 7792
rect 34188 7792 34272 7812
rect 34188 7784 34208 7792
rect 34216 7784 34244 7792
rect 34252 7784 34272 7792
rect 34308 7792 34392 7812
rect 34308 7784 34328 7792
rect 34336 7784 34364 7792
rect 34372 7784 34392 7792
rect 34428 7792 34512 7812
rect 34428 7784 34448 7792
rect 34456 7784 34484 7792
rect 34492 7784 34512 7792
rect 34548 7792 34632 7812
rect 34548 7784 34568 7792
rect 34576 7784 34604 7792
rect 34612 7784 34632 7792
rect 34668 7792 34752 7812
rect 34668 7784 34688 7792
rect 34696 7784 34724 7792
rect 34732 7784 34752 7792
rect 34788 7792 34872 7812
rect 34788 7784 34808 7792
rect 34816 7784 34844 7792
rect 34852 7784 34872 7792
rect 34908 7792 34992 7812
rect 34908 7784 34928 7792
rect 34936 7784 34964 7792
rect 34972 7784 34992 7792
rect 35028 7792 35112 7812
rect 35028 7784 35048 7792
rect 35056 7784 35084 7792
rect 35092 7784 35112 7792
rect 35148 7792 35232 7812
rect 35148 7784 35168 7792
rect 35176 7784 35204 7792
rect 35212 7784 35232 7792
rect 35268 7792 35352 7812
rect 35268 7784 35288 7792
rect 35296 7784 35324 7792
rect 35332 7784 35352 7792
rect 35388 7792 35472 7812
rect 35388 7784 35408 7792
rect 35416 7784 35444 7792
rect 35452 7784 35472 7792
rect 35508 7792 35592 7812
rect 35508 7784 35528 7792
rect 35536 7784 35564 7792
rect 35572 7784 35592 7792
rect 35628 7792 35712 7812
rect 35628 7784 35648 7792
rect 35656 7784 35684 7792
rect 35692 7784 35712 7792
rect 35748 7792 35832 7812
rect 35748 7784 35768 7792
rect 35776 7784 35804 7792
rect 35812 7784 35832 7792
rect 35868 7792 35952 7812
rect 35868 7784 35888 7792
rect 35896 7784 35924 7792
rect 35932 7784 35952 7792
rect 35988 7792 36072 7812
rect 35988 7784 36008 7792
rect 36016 7784 36044 7792
rect 36052 7784 36072 7792
rect 36108 7792 36192 7812
rect 36108 7784 36128 7792
rect 36136 7784 36164 7792
rect 36172 7784 36192 7792
rect 36228 7792 36312 7812
rect 36228 7784 36248 7792
rect 36256 7784 36284 7792
rect 36292 7784 36312 7792
rect 36348 7792 36432 7812
rect 36348 7784 36368 7792
rect 36376 7784 36404 7792
rect 36412 7784 36432 7792
rect 36468 7792 36552 7812
rect 36468 7784 36488 7792
rect 36496 7784 36524 7792
rect 36532 7784 36552 7792
rect 36588 7792 36672 7812
rect 36588 7784 36608 7792
rect 36616 7784 36644 7792
rect 36652 7784 36672 7792
rect 36708 7792 36792 7812
rect 36708 7784 36728 7792
rect 36736 7784 36764 7792
rect 36772 7784 36792 7792
rect 36828 7792 36912 7812
rect 36828 7784 36848 7792
rect 36856 7784 36884 7792
rect 36892 7784 36912 7792
rect 36948 7792 37032 7812
rect 36948 7784 36968 7792
rect 36976 7784 37004 7792
rect 37012 7784 37032 7792
rect 37068 7792 37152 7812
rect 37068 7784 37088 7792
rect 37096 7784 37124 7792
rect 37132 7784 37152 7792
rect 37188 7792 37272 7812
rect 37188 7784 37208 7792
rect 37216 7784 37244 7792
rect 37252 7784 37272 7792
rect 37308 7792 37392 7812
rect 37308 7784 37328 7792
rect 37336 7784 37364 7792
rect 37372 7784 37392 7792
rect 37428 7792 37512 7812
rect 37428 7784 37448 7792
rect 37456 7784 37484 7792
rect 37492 7784 37512 7792
rect 37548 7792 37632 7812
rect 37548 7784 37568 7792
rect 37576 7784 37604 7792
rect 37612 7784 37632 7792
rect 37668 7792 37752 7812
rect 37668 7784 37688 7792
rect 37696 7784 37724 7792
rect 37732 7784 37752 7792
rect 37788 7792 37872 7812
rect 37788 7784 37808 7792
rect 37816 7784 37844 7792
rect 37852 7784 37872 7792
rect 37908 7792 37992 7812
rect 37908 7784 37928 7792
rect 37936 7784 37964 7792
rect 37972 7784 37992 7792
rect 38028 7792 38112 7812
rect 38028 7784 38048 7792
rect 38056 7784 38084 7792
rect 38092 7784 38112 7792
rect 38148 7792 38232 7812
rect 38148 7784 38168 7792
rect 38176 7784 38204 7792
rect 38212 7784 38232 7792
rect 38268 7792 38352 7812
rect 38268 7784 38288 7792
rect 38296 7784 38324 7792
rect 38332 7784 38352 7792
rect 38388 7792 38472 7812
rect 38388 7784 38408 7792
rect 38416 7784 38444 7792
rect 38452 7784 38472 7792
rect 38508 7792 38592 7812
rect 38508 7784 38528 7792
rect 38536 7784 38564 7792
rect 38572 7784 38592 7792
rect 38628 7792 38712 7812
rect 38628 7784 38648 7792
rect 38656 7784 38684 7792
rect 38692 7784 38712 7792
rect 38748 7792 38832 7812
rect 38748 7784 38768 7792
rect 38776 7784 38804 7792
rect 38812 7784 38832 7792
rect 38868 7792 38952 7812
rect 38868 7784 38888 7792
rect 38896 7784 38924 7792
rect 38932 7784 38952 7792
rect 38988 7792 39072 7812
rect 38988 7784 39008 7792
rect 39016 7784 39044 7792
rect 39052 7784 39072 7792
rect 39108 7792 39192 7812
rect 39108 7784 39128 7792
rect 39136 7784 39164 7792
rect 39172 7784 39192 7792
rect 39228 7792 39312 7812
rect 39228 7784 39248 7792
rect 39256 7784 39284 7792
rect 39292 7784 39312 7792
rect 39348 7792 39432 7812
rect 39348 7784 39368 7792
rect 39376 7784 39404 7792
rect 39412 7784 39432 7792
rect 39468 7792 39552 7812
rect 39468 7784 39488 7792
rect 39496 7784 39524 7792
rect 39532 7784 39552 7792
rect 39588 7792 39672 7812
rect 39588 7784 39608 7792
rect 39616 7784 39644 7792
rect 39652 7784 39672 7792
rect 39708 7792 39792 7812
rect 39708 7784 39728 7792
rect 39736 7784 39764 7792
rect 39772 7784 39792 7792
rect 39828 7792 39912 7812
rect 39828 7784 39848 7792
rect 39856 7784 39884 7792
rect 39892 7784 39912 7792
rect 39948 7792 40032 7812
rect 39948 7784 39968 7792
rect 39976 7784 40004 7792
rect 40012 7784 40032 7792
rect 40068 7792 40152 7812
rect 40068 7784 40088 7792
rect 40096 7784 40124 7792
rect 40132 7784 40152 7792
rect 40188 7792 40272 7812
rect 40188 7784 40208 7792
rect 40216 7784 40244 7792
rect 40252 7784 40272 7792
rect 40308 7792 40392 7812
rect 40308 7784 40328 7792
rect 40336 7784 40364 7792
rect 40372 7784 40392 7792
rect 40428 7792 40512 7812
rect 40428 7784 40448 7792
rect 40456 7784 40484 7792
rect 40492 7784 40512 7792
rect 40548 7792 40632 7812
rect 40548 7784 40568 7792
rect 40576 7784 40604 7792
rect 40612 7784 40632 7792
rect 40668 7792 40752 7812
rect 40668 7784 40688 7792
rect 40696 7784 40724 7792
rect 40732 7784 40752 7792
rect 40788 7792 40872 7812
rect 40788 7784 40808 7792
rect 40816 7784 40844 7792
rect 40852 7784 40872 7792
rect 40908 7792 40992 7812
rect 40908 7784 40928 7792
rect 40936 7784 40964 7792
rect 40972 7784 40992 7792
rect 41028 7792 41112 7812
rect 41028 7784 41048 7792
rect 41056 7784 41084 7792
rect 41092 7784 41112 7792
rect 41148 7792 41232 7812
rect 41148 7784 41168 7792
rect 41176 7784 41204 7792
rect 41212 7784 41232 7792
rect 41268 7792 41352 7812
rect 41268 7784 41288 7792
rect 41296 7784 41324 7792
rect 41332 7784 41352 7792
rect 41388 7792 41472 7812
rect 41388 7784 41408 7792
rect 41416 7784 41444 7792
rect 41452 7784 41472 7792
rect 41508 7792 41592 7812
rect 41508 7784 41528 7792
rect 41536 7784 41564 7792
rect 41572 7784 41592 7792
rect 41628 7792 41712 7812
rect 41628 7784 41648 7792
rect 41656 7784 41684 7792
rect 41692 7784 41712 7792
rect 41748 7792 41832 7812
rect 41748 7784 41768 7792
rect 41776 7784 41804 7792
rect 41812 7784 41832 7792
rect 41868 7792 41952 7812
rect 41868 7784 41888 7792
rect 41896 7784 41924 7792
rect 41932 7784 41952 7792
rect 41988 7792 42072 7812
rect 41988 7784 42008 7792
rect 42016 7784 42044 7792
rect 42052 7784 42072 7792
rect 42108 7792 42192 7812
rect 42108 7784 42128 7792
rect 42136 7784 42164 7792
rect 42172 7784 42192 7792
rect 42228 7792 42312 7812
rect 42228 7784 42248 7792
rect 42256 7784 42284 7792
rect 42292 7784 42312 7792
rect 42348 7792 42432 7812
rect 42348 7784 42368 7792
rect 42376 7784 42404 7792
rect 42412 7784 42432 7792
rect 42468 7792 42552 7812
rect 42468 7784 42488 7792
rect 42496 7784 42524 7792
rect 42532 7784 42552 7792
rect 42588 7792 42672 7812
rect 42588 7784 42608 7792
rect 42616 7784 42644 7792
rect 42652 7784 42672 7792
rect 42708 7792 42792 7812
rect 42708 7784 42728 7792
rect 42736 7784 42764 7792
rect 42772 7784 42792 7792
rect 42828 7792 42912 7812
rect 42828 7784 42848 7792
rect 42856 7784 42884 7792
rect 42892 7784 42912 7792
rect 42948 7792 43032 7812
rect 42948 7784 42968 7792
rect 42976 7784 43004 7792
rect 43012 7784 43032 7792
rect 43068 7792 43152 7812
rect 43068 7784 43088 7792
rect 43096 7784 43124 7792
rect 43132 7784 43152 7792
rect 43188 7792 43272 7812
rect 43188 7784 43208 7792
rect 43216 7784 43244 7792
rect 43252 7784 43272 7792
rect 43308 7792 43392 7812
rect 43308 7784 43328 7792
rect 43336 7784 43364 7792
rect 43372 7784 43392 7792
rect 43428 7792 43512 7812
rect 43428 7784 43448 7792
rect 43456 7784 43484 7792
rect 43492 7784 43512 7792
rect 43548 7792 43632 7812
rect 43548 7784 43568 7792
rect 43576 7784 43604 7792
rect 43612 7784 43632 7792
rect 43668 7792 43752 7812
rect 43668 7784 43688 7792
rect 43696 7784 43724 7792
rect 43732 7784 43752 7792
rect 43788 7792 43872 7812
rect 43788 7784 43808 7792
rect 43816 7784 43844 7792
rect 43852 7784 43872 7792
rect 43908 7792 43992 7812
rect 43908 7784 43928 7792
rect 43936 7784 43964 7792
rect 43972 7784 43992 7792
rect 44028 7792 44112 7812
rect 44028 7784 44048 7792
rect 44056 7784 44084 7792
rect 44092 7784 44112 7792
rect 44148 7792 44232 7812
rect 44148 7784 44168 7792
rect 44176 7784 44204 7792
rect 44212 7784 44232 7792
rect 44268 7792 44352 7812
rect 44268 7784 44288 7792
rect 44296 7784 44324 7792
rect 44332 7784 44352 7792
rect 44388 7792 44472 7812
rect 44388 7784 44408 7792
rect 44416 7784 44444 7792
rect 44452 7784 44472 7792
rect 44508 7792 44592 7812
rect 44508 7784 44528 7792
rect 44536 7784 44564 7792
rect 44572 7784 44592 7792
rect 44628 7792 44712 7812
rect 44628 7784 44648 7792
rect 44656 7784 44684 7792
rect 44692 7784 44712 7792
rect 44748 7792 44832 7812
rect 44748 7784 44768 7792
rect 44776 7784 44804 7792
rect 44812 7784 44832 7792
rect 44868 7792 44952 7812
rect 44868 7784 44888 7792
rect 44896 7784 44924 7792
rect 44932 7784 44952 7792
rect 44988 7792 45072 7812
rect 44988 7784 45008 7792
rect 45016 7784 45044 7792
rect 45052 7784 45072 7792
rect 45108 7792 45192 7812
rect 45108 7784 45128 7792
rect 45136 7784 45164 7792
rect 45172 7784 45192 7792
rect 45228 7792 45312 7812
rect 45228 7784 45248 7792
rect 45256 7784 45284 7792
rect 45292 7784 45312 7792
rect 45348 7792 45432 7812
rect 45348 7784 45368 7792
rect 45376 7784 45404 7792
rect 45412 7784 45432 7792
rect 45468 7792 45552 7812
rect 45468 7784 45488 7792
rect 45496 7784 45524 7792
rect 45532 7784 45552 7792
rect 45588 7792 45672 7812
rect 45588 7784 45608 7792
rect 45616 7784 45644 7792
rect 45652 7784 45672 7792
rect 25936 7756 25992 7784
rect 26056 7756 26112 7784
rect 26176 7756 26232 7784
rect 26296 7756 26352 7784
rect 26416 7756 26472 7784
rect 26536 7756 26592 7784
rect 26656 7756 26712 7784
rect 26776 7756 26832 7784
rect 26896 7756 26952 7784
rect 27016 7756 27072 7784
rect 27136 7756 27192 7784
rect 27256 7756 27312 7784
rect 27376 7756 27432 7784
rect 27496 7756 27552 7784
rect 27616 7756 27672 7784
rect 27736 7756 27792 7784
rect 27856 7756 27912 7784
rect 27976 7756 28032 7784
rect 28096 7756 28152 7784
rect 28216 7756 28272 7784
rect 28336 7756 28392 7784
rect 28456 7756 28512 7784
rect 28576 7756 28632 7784
rect 28696 7756 28752 7784
rect 28816 7756 28872 7784
rect 28936 7756 28992 7784
rect 29056 7756 29112 7784
rect 29176 7756 29232 7784
rect 29296 7756 29352 7784
rect 29416 7756 29472 7784
rect 29536 7756 29592 7784
rect 29656 7756 29712 7784
rect 29776 7756 29832 7784
rect 29896 7756 29952 7784
rect 30016 7756 30072 7784
rect 30136 7756 30192 7784
rect 30256 7756 30312 7784
rect 30376 7756 30432 7784
rect 30496 7756 30552 7784
rect 30616 7756 30672 7784
rect 30736 7756 30792 7784
rect 30856 7756 30912 7784
rect 30976 7756 31032 7784
rect 31096 7756 31152 7784
rect 31216 7756 31272 7784
rect 31336 7756 31392 7784
rect 31456 7756 31512 7784
rect 31576 7756 31632 7784
rect 31696 7756 31752 7784
rect 31816 7756 31872 7784
rect 31936 7756 31992 7784
rect 32056 7756 32112 7784
rect 32176 7756 32232 7784
rect 32296 7756 32352 7784
rect 32416 7756 32472 7784
rect 32536 7756 32592 7784
rect 32656 7756 32712 7784
rect 32776 7756 32832 7784
rect 32896 7756 32952 7784
rect 33016 7756 33072 7784
rect 33136 7756 33192 7784
rect 33256 7756 33312 7784
rect 33376 7756 33432 7784
rect 33496 7756 33552 7784
rect 33616 7756 33672 7784
rect 33736 7756 33792 7784
rect 33856 7756 33912 7784
rect 33976 7756 34032 7784
rect 34096 7756 34152 7784
rect 34216 7756 34272 7784
rect 34336 7756 34392 7784
rect 34456 7756 34512 7784
rect 34576 7756 34632 7784
rect 34696 7756 34752 7784
rect 34816 7756 34872 7784
rect 34936 7756 34992 7784
rect 35056 7756 35112 7784
rect 35176 7756 35232 7784
rect 35296 7756 35352 7784
rect 35416 7756 35472 7784
rect 35536 7756 35592 7784
rect 35656 7756 35712 7784
rect 35776 7756 35832 7784
rect 35896 7756 35952 7784
rect 36016 7756 36072 7784
rect 36136 7756 36192 7784
rect 36256 7756 36312 7784
rect 36376 7756 36432 7784
rect 36496 7756 36552 7784
rect 36616 7756 36672 7784
rect 36736 7756 36792 7784
rect 36856 7756 36912 7784
rect 36976 7756 37032 7784
rect 37096 7756 37152 7784
rect 37216 7756 37272 7784
rect 37336 7756 37392 7784
rect 37456 7756 37512 7784
rect 37576 7756 37632 7784
rect 37696 7756 37752 7784
rect 37816 7756 37872 7784
rect 37936 7756 37992 7784
rect 38056 7756 38112 7784
rect 38176 7756 38232 7784
rect 38296 7756 38352 7784
rect 38416 7756 38472 7784
rect 38536 7756 38592 7784
rect 38656 7756 38712 7784
rect 38776 7756 38832 7784
rect 38896 7756 38952 7784
rect 39016 7756 39072 7784
rect 39136 7756 39192 7784
rect 39256 7756 39312 7784
rect 39376 7756 39432 7784
rect 39496 7756 39552 7784
rect 39616 7756 39672 7784
rect 39736 7756 39792 7784
rect 39856 7756 39912 7784
rect 39976 7756 40032 7784
rect 40096 7756 40152 7784
rect 40216 7756 40272 7784
rect 40336 7756 40392 7784
rect 40456 7756 40512 7784
rect 40576 7756 40632 7784
rect 40696 7756 40752 7784
rect 40816 7756 40872 7784
rect 40936 7756 40992 7784
rect 41056 7756 41112 7784
rect 41176 7756 41232 7784
rect 41296 7756 41352 7784
rect 41416 7756 41472 7784
rect 41536 7756 41592 7784
rect 41656 7756 41712 7784
rect 41776 7756 41832 7784
rect 41896 7756 41952 7784
rect 42016 7756 42072 7784
rect 42136 7756 42192 7784
rect 42256 7756 42312 7784
rect 42376 7756 42432 7784
rect 42496 7756 42552 7784
rect 42616 7756 42672 7784
rect 42736 7756 42792 7784
rect 42856 7756 42912 7784
rect 42976 7756 43032 7784
rect 43096 7756 43152 7784
rect 43216 7756 43272 7784
rect 43336 7756 43392 7784
rect 43456 7756 43512 7784
rect 43576 7756 43632 7784
rect 43696 7756 43752 7784
rect 43816 7756 43872 7784
rect 43936 7756 43992 7784
rect 44056 7756 44112 7784
rect 44176 7756 44232 7784
rect 44296 7756 44352 7784
rect 44416 7756 44472 7784
rect 44536 7756 44592 7784
rect 44656 7756 44712 7784
rect 44776 7756 44832 7784
rect 44896 7756 44952 7784
rect 45016 7756 45072 7784
rect 45136 7756 45192 7784
rect 45256 7756 45312 7784
rect 45376 7756 45432 7784
rect 45496 7756 45552 7784
rect 45616 7756 45672 7784
rect 25908 3112 25992 3132
rect 25908 3104 25928 3112
rect 25936 3104 25964 3112
rect 25972 3104 25992 3112
rect 26028 3112 26112 3132
rect 26028 3104 26048 3112
rect 26056 3104 26084 3112
rect 26092 3104 26112 3112
rect 26148 3112 26232 3132
rect 26148 3104 26168 3112
rect 26176 3104 26204 3112
rect 26212 3104 26232 3112
rect 26268 3112 26352 3132
rect 26268 3104 26288 3112
rect 26296 3104 26324 3112
rect 26332 3104 26352 3112
rect 26388 3112 26472 3132
rect 26388 3104 26408 3112
rect 26416 3104 26444 3112
rect 26452 3104 26472 3112
rect 26508 3112 26592 3132
rect 26508 3104 26528 3112
rect 26536 3104 26564 3112
rect 26572 3104 26592 3112
rect 26628 3112 26712 3132
rect 26628 3104 26648 3112
rect 26656 3104 26684 3112
rect 26692 3104 26712 3112
rect 26748 3112 26832 3132
rect 26748 3104 26768 3112
rect 26776 3104 26804 3112
rect 26812 3104 26832 3112
rect 26868 3112 26952 3132
rect 26868 3104 26888 3112
rect 26896 3104 26924 3112
rect 26932 3104 26952 3112
rect 26988 3112 27072 3132
rect 26988 3104 27008 3112
rect 27016 3104 27044 3112
rect 27052 3104 27072 3112
rect 27108 3112 27192 3132
rect 27108 3104 27128 3112
rect 27136 3104 27164 3112
rect 27172 3104 27192 3112
rect 27228 3112 27312 3132
rect 27228 3104 27248 3112
rect 27256 3104 27284 3112
rect 27292 3104 27312 3112
rect 27348 3112 27432 3132
rect 27348 3104 27368 3112
rect 27376 3104 27404 3112
rect 27412 3104 27432 3112
rect 27468 3112 27552 3132
rect 27468 3104 27488 3112
rect 27496 3104 27524 3112
rect 27532 3104 27552 3112
rect 27588 3112 27672 3132
rect 27588 3104 27608 3112
rect 27616 3104 27644 3112
rect 27652 3104 27672 3112
rect 27708 3112 27792 3132
rect 27708 3104 27728 3112
rect 27736 3104 27764 3112
rect 27772 3104 27792 3112
rect 27828 3112 27912 3132
rect 27828 3104 27848 3112
rect 27856 3104 27884 3112
rect 27892 3104 27912 3112
rect 27948 3112 28032 3132
rect 27948 3104 27968 3112
rect 27976 3104 28004 3112
rect 28012 3104 28032 3112
rect 28068 3112 28152 3132
rect 28068 3104 28088 3112
rect 28096 3104 28124 3112
rect 28132 3104 28152 3112
rect 28188 3112 28272 3132
rect 28188 3104 28208 3112
rect 28216 3104 28244 3112
rect 28252 3104 28272 3112
rect 28308 3112 28392 3132
rect 28308 3104 28328 3112
rect 28336 3104 28364 3112
rect 28372 3104 28392 3112
rect 28428 3112 28512 3132
rect 28428 3104 28448 3112
rect 28456 3104 28484 3112
rect 28492 3104 28512 3112
rect 28548 3112 28632 3132
rect 28548 3104 28568 3112
rect 28576 3104 28604 3112
rect 28612 3104 28632 3112
rect 28668 3112 28752 3132
rect 28668 3104 28688 3112
rect 28696 3104 28724 3112
rect 28732 3104 28752 3112
rect 28788 3112 28872 3132
rect 28788 3104 28808 3112
rect 28816 3104 28844 3112
rect 28852 3104 28872 3112
rect 28908 3112 28992 3132
rect 28908 3104 28928 3112
rect 28936 3104 28964 3112
rect 28972 3104 28992 3112
rect 29028 3112 29112 3132
rect 29028 3104 29048 3112
rect 29056 3104 29084 3112
rect 29092 3104 29112 3112
rect 29148 3112 29232 3132
rect 29148 3104 29168 3112
rect 29176 3104 29204 3112
rect 29212 3104 29232 3112
rect 29268 3112 29352 3132
rect 29268 3104 29288 3112
rect 29296 3104 29324 3112
rect 29332 3104 29352 3112
rect 29388 3112 29472 3132
rect 29388 3104 29408 3112
rect 29416 3104 29444 3112
rect 29452 3104 29472 3112
rect 29508 3112 29592 3132
rect 29508 3104 29528 3112
rect 29536 3104 29564 3112
rect 29572 3104 29592 3112
rect 29628 3112 29712 3132
rect 29628 3104 29648 3112
rect 29656 3104 29684 3112
rect 29692 3104 29712 3112
rect 29748 3112 29832 3132
rect 29748 3104 29768 3112
rect 29776 3104 29804 3112
rect 29812 3104 29832 3112
rect 29868 3112 29952 3132
rect 29868 3104 29888 3112
rect 29896 3104 29924 3112
rect 29932 3104 29952 3112
rect 29988 3112 30072 3132
rect 29988 3104 30008 3112
rect 30016 3104 30044 3112
rect 30052 3104 30072 3112
rect 30108 3112 30192 3132
rect 30108 3104 30128 3112
rect 30136 3104 30164 3112
rect 30172 3104 30192 3112
rect 30228 3112 30312 3132
rect 30228 3104 30248 3112
rect 30256 3104 30284 3112
rect 30292 3104 30312 3112
rect 30348 3112 30432 3132
rect 30348 3104 30368 3112
rect 30376 3104 30404 3112
rect 30412 3104 30432 3112
rect 30468 3112 30552 3132
rect 30468 3104 30488 3112
rect 30496 3104 30524 3112
rect 30532 3104 30552 3112
rect 30588 3112 30672 3132
rect 30588 3104 30608 3112
rect 30616 3104 30644 3112
rect 30652 3104 30672 3112
rect 30708 3112 30792 3132
rect 30708 3104 30728 3112
rect 30736 3104 30764 3112
rect 30772 3104 30792 3112
rect 30828 3112 30912 3132
rect 30828 3104 30848 3112
rect 30856 3104 30884 3112
rect 30892 3104 30912 3112
rect 30948 3112 31032 3132
rect 30948 3104 30968 3112
rect 30976 3104 31004 3112
rect 31012 3104 31032 3112
rect 31068 3112 31152 3132
rect 31068 3104 31088 3112
rect 31096 3104 31124 3112
rect 31132 3104 31152 3112
rect 31188 3112 31272 3132
rect 31188 3104 31208 3112
rect 31216 3104 31244 3112
rect 31252 3104 31272 3112
rect 31308 3112 31392 3132
rect 31308 3104 31328 3112
rect 31336 3104 31364 3112
rect 31372 3104 31392 3112
rect 31428 3112 31512 3132
rect 31428 3104 31448 3112
rect 31456 3104 31484 3112
rect 31492 3104 31512 3112
rect 31548 3112 31632 3132
rect 31548 3104 31568 3112
rect 31576 3104 31604 3112
rect 31612 3104 31632 3112
rect 31668 3112 31752 3132
rect 31668 3104 31688 3112
rect 31696 3104 31724 3112
rect 31732 3104 31752 3112
rect 31788 3112 31872 3132
rect 31788 3104 31808 3112
rect 31816 3104 31844 3112
rect 31852 3104 31872 3112
rect 31908 3112 31992 3132
rect 31908 3104 31928 3112
rect 31936 3104 31964 3112
rect 31972 3104 31992 3112
rect 32028 3112 32112 3132
rect 32028 3104 32048 3112
rect 32056 3104 32084 3112
rect 32092 3104 32112 3112
rect 32148 3112 32232 3132
rect 32148 3104 32168 3112
rect 32176 3104 32204 3112
rect 32212 3104 32232 3112
rect 32268 3112 32352 3132
rect 32268 3104 32288 3112
rect 32296 3104 32324 3112
rect 32332 3104 32352 3112
rect 32388 3112 32472 3132
rect 32388 3104 32408 3112
rect 32416 3104 32444 3112
rect 32452 3104 32472 3112
rect 32508 3112 32592 3132
rect 32508 3104 32528 3112
rect 32536 3104 32564 3112
rect 32572 3104 32592 3112
rect 32628 3112 32712 3132
rect 32628 3104 32648 3112
rect 32656 3104 32684 3112
rect 32692 3104 32712 3112
rect 32748 3112 32832 3132
rect 32748 3104 32768 3112
rect 32776 3104 32804 3112
rect 32812 3104 32832 3112
rect 32868 3112 32952 3132
rect 32868 3104 32888 3112
rect 32896 3104 32924 3112
rect 32932 3104 32952 3112
rect 32988 3112 33072 3132
rect 32988 3104 33008 3112
rect 33016 3104 33044 3112
rect 33052 3104 33072 3112
rect 33108 3112 33192 3132
rect 33108 3104 33128 3112
rect 33136 3104 33164 3112
rect 33172 3104 33192 3112
rect 33228 3112 33312 3132
rect 33228 3104 33248 3112
rect 33256 3104 33284 3112
rect 33292 3104 33312 3112
rect 33348 3112 33432 3132
rect 33348 3104 33368 3112
rect 33376 3104 33404 3112
rect 33412 3104 33432 3112
rect 33468 3112 33552 3132
rect 33468 3104 33488 3112
rect 33496 3104 33524 3112
rect 33532 3104 33552 3112
rect 33588 3112 33672 3132
rect 33588 3104 33608 3112
rect 33616 3104 33644 3112
rect 33652 3104 33672 3112
rect 33708 3112 33792 3132
rect 33708 3104 33728 3112
rect 33736 3104 33764 3112
rect 33772 3104 33792 3112
rect 33828 3112 33912 3132
rect 33828 3104 33848 3112
rect 33856 3104 33884 3112
rect 33892 3104 33912 3112
rect 33948 3112 34032 3132
rect 33948 3104 33968 3112
rect 33976 3104 34004 3112
rect 34012 3104 34032 3112
rect 34068 3112 34152 3132
rect 34068 3104 34088 3112
rect 34096 3104 34124 3112
rect 34132 3104 34152 3112
rect 34188 3112 34272 3132
rect 34188 3104 34208 3112
rect 34216 3104 34244 3112
rect 34252 3104 34272 3112
rect 34308 3112 34392 3132
rect 34308 3104 34328 3112
rect 34336 3104 34364 3112
rect 34372 3104 34392 3112
rect 34428 3112 34512 3132
rect 34428 3104 34448 3112
rect 34456 3104 34484 3112
rect 34492 3104 34512 3112
rect 34548 3112 34632 3132
rect 34548 3104 34568 3112
rect 34576 3104 34604 3112
rect 34612 3104 34632 3112
rect 34668 3112 34752 3132
rect 34668 3104 34688 3112
rect 34696 3104 34724 3112
rect 34732 3104 34752 3112
rect 34788 3112 34872 3132
rect 34788 3104 34808 3112
rect 34816 3104 34844 3112
rect 34852 3104 34872 3112
rect 34908 3112 34992 3132
rect 34908 3104 34928 3112
rect 34936 3104 34964 3112
rect 34972 3104 34992 3112
rect 35028 3112 35112 3132
rect 35028 3104 35048 3112
rect 35056 3104 35084 3112
rect 35092 3104 35112 3112
rect 35148 3112 35232 3132
rect 35148 3104 35168 3112
rect 35176 3104 35204 3112
rect 35212 3104 35232 3112
rect 35268 3112 35352 3132
rect 35268 3104 35288 3112
rect 35296 3104 35324 3112
rect 35332 3104 35352 3112
rect 35388 3112 35472 3132
rect 35388 3104 35408 3112
rect 35416 3104 35444 3112
rect 35452 3104 35472 3112
rect 35508 3112 35592 3132
rect 35508 3104 35528 3112
rect 35536 3104 35564 3112
rect 35572 3104 35592 3112
rect 35628 3112 35712 3132
rect 35628 3104 35648 3112
rect 35656 3104 35684 3112
rect 35692 3104 35712 3112
rect 35748 3112 35832 3132
rect 35748 3104 35768 3112
rect 35776 3104 35804 3112
rect 35812 3104 35832 3112
rect 35868 3112 35952 3132
rect 35868 3104 35888 3112
rect 35896 3104 35924 3112
rect 35932 3104 35952 3112
rect 35988 3112 36072 3132
rect 35988 3104 36008 3112
rect 36016 3104 36044 3112
rect 36052 3104 36072 3112
rect 36108 3112 36192 3132
rect 36108 3104 36128 3112
rect 36136 3104 36164 3112
rect 36172 3104 36192 3112
rect 36228 3112 36312 3132
rect 36228 3104 36248 3112
rect 36256 3104 36284 3112
rect 36292 3104 36312 3112
rect 36348 3112 36432 3132
rect 36348 3104 36368 3112
rect 36376 3104 36404 3112
rect 36412 3104 36432 3112
rect 36468 3112 36552 3132
rect 36468 3104 36488 3112
rect 36496 3104 36524 3112
rect 36532 3104 36552 3112
rect 36588 3112 36672 3132
rect 36588 3104 36608 3112
rect 36616 3104 36644 3112
rect 36652 3104 36672 3112
rect 36708 3112 36792 3132
rect 36708 3104 36728 3112
rect 36736 3104 36764 3112
rect 36772 3104 36792 3112
rect 36828 3112 36912 3132
rect 36828 3104 36848 3112
rect 36856 3104 36884 3112
rect 36892 3104 36912 3112
rect 36948 3112 37032 3132
rect 36948 3104 36968 3112
rect 36976 3104 37004 3112
rect 37012 3104 37032 3112
rect 37068 3112 37152 3132
rect 37068 3104 37088 3112
rect 37096 3104 37124 3112
rect 37132 3104 37152 3112
rect 37188 3112 37272 3132
rect 37188 3104 37208 3112
rect 37216 3104 37244 3112
rect 37252 3104 37272 3112
rect 37308 3112 37392 3132
rect 37308 3104 37328 3112
rect 37336 3104 37364 3112
rect 37372 3104 37392 3112
rect 37428 3112 37512 3132
rect 37428 3104 37448 3112
rect 37456 3104 37484 3112
rect 37492 3104 37512 3112
rect 37548 3112 37632 3132
rect 37548 3104 37568 3112
rect 37576 3104 37604 3112
rect 37612 3104 37632 3112
rect 37668 3112 37752 3132
rect 37668 3104 37688 3112
rect 37696 3104 37724 3112
rect 37732 3104 37752 3112
rect 37788 3112 37872 3132
rect 37788 3104 37808 3112
rect 37816 3104 37844 3112
rect 37852 3104 37872 3112
rect 37908 3112 37992 3132
rect 37908 3104 37928 3112
rect 37936 3104 37964 3112
rect 37972 3104 37992 3112
rect 38028 3112 38112 3132
rect 38028 3104 38048 3112
rect 38056 3104 38084 3112
rect 38092 3104 38112 3112
rect 38148 3112 38232 3132
rect 38148 3104 38168 3112
rect 38176 3104 38204 3112
rect 38212 3104 38232 3112
rect 38268 3112 38352 3132
rect 38268 3104 38288 3112
rect 38296 3104 38324 3112
rect 38332 3104 38352 3112
rect 38388 3112 38472 3132
rect 38388 3104 38408 3112
rect 38416 3104 38444 3112
rect 38452 3104 38472 3112
rect 38508 3112 38592 3132
rect 38508 3104 38528 3112
rect 38536 3104 38564 3112
rect 38572 3104 38592 3112
rect 38628 3112 38712 3132
rect 38628 3104 38648 3112
rect 38656 3104 38684 3112
rect 38692 3104 38712 3112
rect 38748 3112 38832 3132
rect 38748 3104 38768 3112
rect 38776 3104 38804 3112
rect 38812 3104 38832 3112
rect 38868 3112 38952 3132
rect 38868 3104 38888 3112
rect 38896 3104 38924 3112
rect 38932 3104 38952 3112
rect 38988 3112 39072 3132
rect 38988 3104 39008 3112
rect 39016 3104 39044 3112
rect 39052 3104 39072 3112
rect 39108 3112 39192 3132
rect 39108 3104 39128 3112
rect 39136 3104 39164 3112
rect 39172 3104 39192 3112
rect 39228 3112 39312 3132
rect 39228 3104 39248 3112
rect 39256 3104 39284 3112
rect 39292 3104 39312 3112
rect 39348 3112 39432 3132
rect 39348 3104 39368 3112
rect 39376 3104 39404 3112
rect 39412 3104 39432 3112
rect 39468 3112 39552 3132
rect 39468 3104 39488 3112
rect 39496 3104 39524 3112
rect 39532 3104 39552 3112
rect 39588 3112 39672 3132
rect 39588 3104 39608 3112
rect 39616 3104 39644 3112
rect 39652 3104 39672 3112
rect 39708 3112 39792 3132
rect 39708 3104 39728 3112
rect 39736 3104 39764 3112
rect 39772 3104 39792 3112
rect 39828 3112 39912 3132
rect 39828 3104 39848 3112
rect 39856 3104 39884 3112
rect 39892 3104 39912 3112
rect 39948 3112 40032 3132
rect 39948 3104 39968 3112
rect 39976 3104 40004 3112
rect 40012 3104 40032 3112
rect 40068 3112 40152 3132
rect 40068 3104 40088 3112
rect 40096 3104 40124 3112
rect 40132 3104 40152 3112
rect 40188 3112 40272 3132
rect 40188 3104 40208 3112
rect 40216 3104 40244 3112
rect 40252 3104 40272 3112
rect 40308 3112 40392 3132
rect 40308 3104 40328 3112
rect 40336 3104 40364 3112
rect 40372 3104 40392 3112
rect 40428 3112 40512 3132
rect 40428 3104 40448 3112
rect 40456 3104 40484 3112
rect 40492 3104 40512 3112
rect 40548 3112 40632 3132
rect 40548 3104 40568 3112
rect 40576 3104 40604 3112
rect 40612 3104 40632 3112
rect 40668 3112 40752 3132
rect 40668 3104 40688 3112
rect 40696 3104 40724 3112
rect 40732 3104 40752 3112
rect 40788 3112 40872 3132
rect 40788 3104 40808 3112
rect 40816 3104 40844 3112
rect 40852 3104 40872 3112
rect 40908 3112 40992 3132
rect 40908 3104 40928 3112
rect 40936 3104 40964 3112
rect 40972 3104 40992 3112
rect 41028 3112 41112 3132
rect 41028 3104 41048 3112
rect 41056 3104 41084 3112
rect 41092 3104 41112 3112
rect 41148 3112 41232 3132
rect 41148 3104 41168 3112
rect 41176 3104 41204 3112
rect 41212 3104 41232 3112
rect 41268 3112 41352 3132
rect 41268 3104 41288 3112
rect 41296 3104 41324 3112
rect 41332 3104 41352 3112
rect 41388 3112 41472 3132
rect 41388 3104 41408 3112
rect 41416 3104 41444 3112
rect 41452 3104 41472 3112
rect 41508 3112 41592 3132
rect 41508 3104 41528 3112
rect 41536 3104 41564 3112
rect 41572 3104 41592 3112
rect 41628 3112 41712 3132
rect 41628 3104 41648 3112
rect 41656 3104 41684 3112
rect 41692 3104 41712 3112
rect 41748 3112 41832 3132
rect 41748 3104 41768 3112
rect 41776 3104 41804 3112
rect 41812 3104 41832 3112
rect 41868 3112 41952 3132
rect 41868 3104 41888 3112
rect 41896 3104 41924 3112
rect 41932 3104 41952 3112
rect 41988 3112 42072 3132
rect 41988 3104 42008 3112
rect 42016 3104 42044 3112
rect 42052 3104 42072 3112
rect 42108 3112 42192 3132
rect 42108 3104 42128 3112
rect 42136 3104 42164 3112
rect 42172 3104 42192 3112
rect 42228 3112 42312 3132
rect 42228 3104 42248 3112
rect 42256 3104 42284 3112
rect 42292 3104 42312 3112
rect 42348 3112 42432 3132
rect 42348 3104 42368 3112
rect 42376 3104 42404 3112
rect 42412 3104 42432 3112
rect 42468 3112 42552 3132
rect 42468 3104 42488 3112
rect 42496 3104 42524 3112
rect 42532 3104 42552 3112
rect 42588 3112 42672 3132
rect 42588 3104 42608 3112
rect 42616 3104 42644 3112
rect 42652 3104 42672 3112
rect 42708 3112 42792 3132
rect 42708 3104 42728 3112
rect 42736 3104 42764 3112
rect 42772 3104 42792 3112
rect 42828 3112 42912 3132
rect 42828 3104 42848 3112
rect 42856 3104 42884 3112
rect 42892 3104 42912 3112
rect 42948 3112 43032 3132
rect 42948 3104 42968 3112
rect 42976 3104 43004 3112
rect 43012 3104 43032 3112
rect 43068 3112 43152 3132
rect 43068 3104 43088 3112
rect 43096 3104 43124 3112
rect 43132 3104 43152 3112
rect 43188 3112 43272 3132
rect 43188 3104 43208 3112
rect 43216 3104 43244 3112
rect 43252 3104 43272 3112
rect 43308 3112 43392 3132
rect 43308 3104 43328 3112
rect 43336 3104 43364 3112
rect 43372 3104 43392 3112
rect 43428 3112 43512 3132
rect 43428 3104 43448 3112
rect 43456 3104 43484 3112
rect 43492 3104 43512 3112
rect 43548 3112 43632 3132
rect 43548 3104 43568 3112
rect 43576 3104 43604 3112
rect 43612 3104 43632 3112
rect 43668 3112 43752 3132
rect 43668 3104 43688 3112
rect 43696 3104 43724 3112
rect 43732 3104 43752 3112
rect 43788 3112 43872 3132
rect 43788 3104 43808 3112
rect 43816 3104 43844 3112
rect 43852 3104 43872 3112
rect 43908 3112 43992 3132
rect 43908 3104 43928 3112
rect 43936 3104 43964 3112
rect 43972 3104 43992 3112
rect 44028 3112 44112 3132
rect 44028 3104 44048 3112
rect 44056 3104 44084 3112
rect 44092 3104 44112 3112
rect 44148 3112 44232 3132
rect 44148 3104 44168 3112
rect 44176 3104 44204 3112
rect 44212 3104 44232 3112
rect 44268 3112 44352 3132
rect 44268 3104 44288 3112
rect 44296 3104 44324 3112
rect 44332 3104 44352 3112
rect 44388 3112 44472 3132
rect 44388 3104 44408 3112
rect 44416 3104 44444 3112
rect 44452 3104 44472 3112
rect 44508 3112 44592 3132
rect 44508 3104 44528 3112
rect 44536 3104 44564 3112
rect 44572 3104 44592 3112
rect 44628 3112 44712 3132
rect 44628 3104 44648 3112
rect 44656 3104 44684 3112
rect 44692 3104 44712 3112
rect 44748 3112 44832 3132
rect 44748 3104 44768 3112
rect 44776 3104 44804 3112
rect 44812 3104 44832 3112
rect 44868 3112 44952 3132
rect 44868 3104 44888 3112
rect 44896 3104 44924 3112
rect 44932 3104 44952 3112
rect 44988 3112 45072 3132
rect 44988 3104 45008 3112
rect 45016 3104 45044 3112
rect 45052 3104 45072 3112
rect 45108 3112 45192 3132
rect 45108 3104 45128 3112
rect 45136 3104 45164 3112
rect 45172 3104 45192 3112
rect 45228 3112 45312 3132
rect 45228 3104 45248 3112
rect 45256 3104 45284 3112
rect 45292 3104 45312 3112
rect 45348 3112 45432 3132
rect 45348 3104 45368 3112
rect 45376 3104 45404 3112
rect 45412 3104 45432 3112
rect 45468 3112 45552 3132
rect 45468 3104 45488 3112
rect 45496 3104 45524 3112
rect 45532 3104 45552 3112
rect 45588 3112 45672 3132
rect 45588 3104 45608 3112
rect 45616 3104 45644 3112
rect 45652 3104 45672 3112
rect 25936 3076 25992 3104
rect 26056 3076 26112 3104
rect 26176 3076 26232 3104
rect 26296 3076 26352 3104
rect 26416 3076 26472 3104
rect 26536 3076 26592 3104
rect 26656 3076 26712 3104
rect 26776 3076 26832 3104
rect 26896 3076 26952 3104
rect 27016 3076 27072 3104
rect 27136 3076 27192 3104
rect 27256 3076 27312 3104
rect 27376 3076 27432 3104
rect 27496 3076 27552 3104
rect 27616 3076 27672 3104
rect 27736 3076 27792 3104
rect 27856 3076 27912 3104
rect 27976 3076 28032 3104
rect 28096 3076 28152 3104
rect 28216 3076 28272 3104
rect 28336 3076 28392 3104
rect 28456 3076 28512 3104
rect 28576 3076 28632 3104
rect 28696 3076 28752 3104
rect 28816 3076 28872 3104
rect 28936 3076 28992 3104
rect 29056 3076 29112 3104
rect 29176 3076 29232 3104
rect 29296 3076 29352 3104
rect 29416 3076 29472 3104
rect 29536 3076 29592 3104
rect 29656 3076 29712 3104
rect 29776 3076 29832 3104
rect 29896 3076 29952 3104
rect 30016 3076 30072 3104
rect 30136 3076 30192 3104
rect 30256 3076 30312 3104
rect 30376 3076 30432 3104
rect 30496 3076 30552 3104
rect 30616 3076 30672 3104
rect 30736 3076 30792 3104
rect 30856 3076 30912 3104
rect 30976 3076 31032 3104
rect 31096 3076 31152 3104
rect 31216 3076 31272 3104
rect 31336 3076 31392 3104
rect 31456 3076 31512 3104
rect 31576 3076 31632 3104
rect 31696 3076 31752 3104
rect 31816 3076 31872 3104
rect 31936 3076 31992 3104
rect 32056 3076 32112 3104
rect 32176 3076 32232 3104
rect 32296 3076 32352 3104
rect 32416 3076 32472 3104
rect 32536 3076 32592 3104
rect 32656 3076 32712 3104
rect 32776 3076 32832 3104
rect 32896 3076 32952 3104
rect 33016 3076 33072 3104
rect 33136 3076 33192 3104
rect 33256 3076 33312 3104
rect 33376 3076 33432 3104
rect 33496 3076 33552 3104
rect 33616 3076 33672 3104
rect 33736 3076 33792 3104
rect 33856 3076 33912 3104
rect 33976 3076 34032 3104
rect 34096 3076 34152 3104
rect 34216 3076 34272 3104
rect 34336 3076 34392 3104
rect 34456 3076 34512 3104
rect 34576 3076 34632 3104
rect 34696 3076 34752 3104
rect 34816 3076 34872 3104
rect 34936 3076 34992 3104
rect 35056 3076 35112 3104
rect 35176 3076 35232 3104
rect 35296 3076 35352 3104
rect 35416 3076 35472 3104
rect 35536 3076 35592 3104
rect 35656 3076 35712 3104
rect 35776 3076 35832 3104
rect 35896 3076 35952 3104
rect 36016 3076 36072 3104
rect 36136 3076 36192 3104
rect 36256 3076 36312 3104
rect 36376 3076 36432 3104
rect 36496 3076 36552 3104
rect 36616 3076 36672 3104
rect 36736 3076 36792 3104
rect 36856 3076 36912 3104
rect 36976 3076 37032 3104
rect 37096 3076 37152 3104
rect 37216 3076 37272 3104
rect 37336 3076 37392 3104
rect 37456 3076 37512 3104
rect 37576 3076 37632 3104
rect 37696 3076 37752 3104
rect 37816 3076 37872 3104
rect 37936 3076 37992 3104
rect 38056 3076 38112 3104
rect 38176 3076 38232 3104
rect 38296 3076 38352 3104
rect 38416 3076 38472 3104
rect 38536 3076 38592 3104
rect 38656 3076 38712 3104
rect 38776 3076 38832 3104
rect 38896 3076 38952 3104
rect 39016 3076 39072 3104
rect 39136 3076 39192 3104
rect 39256 3076 39312 3104
rect 39376 3076 39432 3104
rect 39496 3076 39552 3104
rect 39616 3076 39672 3104
rect 39736 3076 39792 3104
rect 39856 3076 39912 3104
rect 39976 3076 40032 3104
rect 40096 3076 40152 3104
rect 40216 3076 40272 3104
rect 40336 3076 40392 3104
rect 40456 3076 40512 3104
rect 40576 3076 40632 3104
rect 40696 3076 40752 3104
rect 40816 3076 40872 3104
rect 40936 3076 40992 3104
rect 41056 3076 41112 3104
rect 41176 3076 41232 3104
rect 41296 3076 41352 3104
rect 41416 3076 41472 3104
rect 41536 3076 41592 3104
rect 41656 3076 41712 3104
rect 41776 3076 41832 3104
rect 41896 3076 41952 3104
rect 42016 3076 42072 3104
rect 42136 3076 42192 3104
rect 42256 3076 42312 3104
rect 42376 3076 42432 3104
rect 42496 3076 42552 3104
rect 42616 3076 42672 3104
rect 42736 3076 42792 3104
rect 42856 3076 42912 3104
rect 42976 3076 43032 3104
rect 43096 3076 43152 3104
rect 43216 3076 43272 3104
rect 43336 3076 43392 3104
rect 43456 3076 43512 3104
rect 43576 3076 43632 3104
rect 43696 3076 43752 3104
rect 43816 3076 43872 3104
rect 43936 3076 43992 3104
rect 44056 3076 44112 3104
rect 44176 3076 44232 3104
rect 44296 3076 44352 3104
rect 44416 3076 44472 3104
rect 44536 3076 44592 3104
rect 44656 3076 44712 3104
rect 44776 3076 44832 3104
rect 44896 3076 44952 3104
rect 45016 3076 45072 3104
rect 45136 3076 45192 3104
rect 45256 3076 45312 3104
rect 45376 3076 45432 3104
rect 45496 3076 45552 3104
rect 45616 3076 45672 3104
rect 25908 2932 25992 2952
rect 25908 2924 25928 2932
rect 25936 2924 25964 2932
rect 25972 2924 25992 2932
rect 26028 2932 26112 2952
rect 26028 2924 26048 2932
rect 26056 2924 26084 2932
rect 26092 2924 26112 2932
rect 26148 2932 26232 2952
rect 26148 2924 26168 2932
rect 26176 2924 26204 2932
rect 26212 2924 26232 2932
rect 26268 2932 26352 2952
rect 26268 2924 26288 2932
rect 26296 2924 26324 2932
rect 26332 2924 26352 2932
rect 26388 2932 26472 2952
rect 26388 2924 26408 2932
rect 26416 2924 26444 2932
rect 26452 2924 26472 2932
rect 26508 2932 26592 2952
rect 26508 2924 26528 2932
rect 26536 2924 26564 2932
rect 26572 2924 26592 2932
rect 26628 2932 26712 2952
rect 26628 2924 26648 2932
rect 26656 2924 26684 2932
rect 26692 2924 26712 2932
rect 26748 2932 26832 2952
rect 26748 2924 26768 2932
rect 26776 2924 26804 2932
rect 26812 2924 26832 2932
rect 26868 2932 26952 2952
rect 26868 2924 26888 2932
rect 26896 2924 26924 2932
rect 26932 2924 26952 2932
rect 26988 2932 27072 2952
rect 26988 2924 27008 2932
rect 27016 2924 27044 2932
rect 27052 2924 27072 2932
rect 27108 2932 27192 2952
rect 27108 2924 27128 2932
rect 27136 2924 27164 2932
rect 27172 2924 27192 2932
rect 27228 2932 27312 2952
rect 27228 2924 27248 2932
rect 27256 2924 27284 2932
rect 27292 2924 27312 2932
rect 27348 2932 27432 2952
rect 27348 2924 27368 2932
rect 27376 2924 27404 2932
rect 27412 2924 27432 2932
rect 27468 2932 27552 2952
rect 27468 2924 27488 2932
rect 27496 2924 27524 2932
rect 27532 2924 27552 2932
rect 27588 2932 27672 2952
rect 27588 2924 27608 2932
rect 27616 2924 27644 2932
rect 27652 2924 27672 2932
rect 27708 2932 27792 2952
rect 27708 2924 27728 2932
rect 27736 2924 27764 2932
rect 27772 2924 27792 2932
rect 27828 2932 27912 2952
rect 27828 2924 27848 2932
rect 27856 2924 27884 2932
rect 27892 2924 27912 2932
rect 27948 2932 28032 2952
rect 27948 2924 27968 2932
rect 27976 2924 28004 2932
rect 28012 2924 28032 2932
rect 28068 2932 28152 2952
rect 28068 2924 28088 2932
rect 28096 2924 28124 2932
rect 28132 2924 28152 2932
rect 28188 2932 28272 2952
rect 28188 2924 28208 2932
rect 28216 2924 28244 2932
rect 28252 2924 28272 2932
rect 28308 2932 28392 2952
rect 28308 2924 28328 2932
rect 28336 2924 28364 2932
rect 28372 2924 28392 2932
rect 28428 2932 28512 2952
rect 28428 2924 28448 2932
rect 28456 2924 28484 2932
rect 28492 2924 28512 2932
rect 28548 2932 28632 2952
rect 28548 2924 28568 2932
rect 28576 2924 28604 2932
rect 28612 2924 28632 2932
rect 28668 2932 28752 2952
rect 28668 2924 28688 2932
rect 28696 2924 28724 2932
rect 28732 2924 28752 2932
rect 28788 2932 28872 2952
rect 28788 2924 28808 2932
rect 28816 2924 28844 2932
rect 28852 2924 28872 2932
rect 28908 2932 28992 2952
rect 28908 2924 28928 2932
rect 28936 2924 28964 2932
rect 28972 2924 28992 2932
rect 29028 2932 29112 2952
rect 29028 2924 29048 2932
rect 29056 2924 29084 2932
rect 29092 2924 29112 2932
rect 29148 2932 29232 2952
rect 29148 2924 29168 2932
rect 29176 2924 29204 2932
rect 29212 2924 29232 2932
rect 29268 2932 29352 2952
rect 29268 2924 29288 2932
rect 29296 2924 29324 2932
rect 29332 2924 29352 2932
rect 29388 2932 29472 2952
rect 29388 2924 29408 2932
rect 29416 2924 29444 2932
rect 29452 2924 29472 2932
rect 29508 2932 29592 2952
rect 29508 2924 29528 2932
rect 29536 2924 29564 2932
rect 29572 2924 29592 2932
rect 29628 2932 29712 2952
rect 29628 2924 29648 2932
rect 29656 2924 29684 2932
rect 29692 2924 29712 2932
rect 29748 2932 29832 2952
rect 29748 2924 29768 2932
rect 29776 2924 29804 2932
rect 29812 2924 29832 2932
rect 29868 2932 29952 2952
rect 29868 2924 29888 2932
rect 29896 2924 29924 2932
rect 29932 2924 29952 2932
rect 29988 2932 30072 2952
rect 29988 2924 30008 2932
rect 30016 2924 30044 2932
rect 30052 2924 30072 2932
rect 30108 2932 30192 2952
rect 30108 2924 30128 2932
rect 30136 2924 30164 2932
rect 30172 2924 30192 2932
rect 30228 2932 30312 2952
rect 30228 2924 30248 2932
rect 30256 2924 30284 2932
rect 30292 2924 30312 2932
rect 30348 2932 30432 2952
rect 30348 2924 30368 2932
rect 30376 2924 30404 2932
rect 30412 2924 30432 2932
rect 30468 2932 30552 2952
rect 30468 2924 30488 2932
rect 30496 2924 30524 2932
rect 30532 2924 30552 2932
rect 30588 2932 30672 2952
rect 30588 2924 30608 2932
rect 30616 2924 30644 2932
rect 30652 2924 30672 2932
rect 30708 2932 30792 2952
rect 30708 2924 30728 2932
rect 30736 2924 30764 2932
rect 30772 2924 30792 2932
rect 30828 2932 30912 2952
rect 30828 2924 30848 2932
rect 30856 2924 30884 2932
rect 30892 2924 30912 2932
rect 30948 2932 31032 2952
rect 30948 2924 30968 2932
rect 30976 2924 31004 2932
rect 31012 2924 31032 2932
rect 31068 2932 31152 2952
rect 31068 2924 31088 2932
rect 31096 2924 31124 2932
rect 31132 2924 31152 2932
rect 31188 2932 31272 2952
rect 31188 2924 31208 2932
rect 31216 2924 31244 2932
rect 31252 2924 31272 2932
rect 31308 2932 31392 2952
rect 31308 2924 31328 2932
rect 31336 2924 31364 2932
rect 31372 2924 31392 2932
rect 31428 2932 31512 2952
rect 31428 2924 31448 2932
rect 31456 2924 31484 2932
rect 31492 2924 31512 2932
rect 31548 2932 31632 2952
rect 31548 2924 31568 2932
rect 31576 2924 31604 2932
rect 31612 2924 31632 2932
rect 31668 2932 31752 2952
rect 31668 2924 31688 2932
rect 31696 2924 31724 2932
rect 31732 2924 31752 2932
rect 31788 2932 31872 2952
rect 31788 2924 31808 2932
rect 31816 2924 31844 2932
rect 31852 2924 31872 2932
rect 31908 2932 31992 2952
rect 31908 2924 31928 2932
rect 31936 2924 31964 2932
rect 31972 2924 31992 2932
rect 32028 2932 32112 2952
rect 32028 2924 32048 2932
rect 32056 2924 32084 2932
rect 32092 2924 32112 2932
rect 32148 2932 32232 2952
rect 32148 2924 32168 2932
rect 32176 2924 32204 2932
rect 32212 2924 32232 2932
rect 32268 2932 32352 2952
rect 32268 2924 32288 2932
rect 32296 2924 32324 2932
rect 32332 2924 32352 2932
rect 32388 2932 32472 2952
rect 32388 2924 32408 2932
rect 32416 2924 32444 2932
rect 32452 2924 32472 2932
rect 32508 2932 32592 2952
rect 32508 2924 32528 2932
rect 32536 2924 32564 2932
rect 32572 2924 32592 2932
rect 32628 2932 32712 2952
rect 32628 2924 32648 2932
rect 32656 2924 32684 2932
rect 32692 2924 32712 2932
rect 32748 2932 32832 2952
rect 32748 2924 32768 2932
rect 32776 2924 32804 2932
rect 32812 2924 32832 2932
rect 32868 2932 32952 2952
rect 32868 2924 32888 2932
rect 32896 2924 32924 2932
rect 32932 2924 32952 2932
rect 32988 2932 33072 2952
rect 32988 2924 33008 2932
rect 33016 2924 33044 2932
rect 33052 2924 33072 2932
rect 33108 2932 33192 2952
rect 33108 2924 33128 2932
rect 33136 2924 33164 2932
rect 33172 2924 33192 2932
rect 33228 2932 33312 2952
rect 33228 2924 33248 2932
rect 33256 2924 33284 2932
rect 33292 2924 33312 2932
rect 33348 2932 33432 2952
rect 33348 2924 33368 2932
rect 33376 2924 33404 2932
rect 33412 2924 33432 2932
rect 33468 2932 33552 2952
rect 33468 2924 33488 2932
rect 33496 2924 33524 2932
rect 33532 2924 33552 2932
rect 33588 2932 33672 2952
rect 33588 2924 33608 2932
rect 33616 2924 33644 2932
rect 33652 2924 33672 2932
rect 33708 2932 33792 2952
rect 33708 2924 33728 2932
rect 33736 2924 33764 2932
rect 33772 2924 33792 2932
rect 33828 2932 33912 2952
rect 33828 2924 33848 2932
rect 33856 2924 33884 2932
rect 33892 2924 33912 2932
rect 33948 2932 34032 2952
rect 33948 2924 33968 2932
rect 33976 2924 34004 2932
rect 34012 2924 34032 2932
rect 34068 2932 34152 2952
rect 34068 2924 34088 2932
rect 34096 2924 34124 2932
rect 34132 2924 34152 2932
rect 34188 2932 34272 2952
rect 34188 2924 34208 2932
rect 34216 2924 34244 2932
rect 34252 2924 34272 2932
rect 34308 2932 34392 2952
rect 34308 2924 34328 2932
rect 34336 2924 34364 2932
rect 34372 2924 34392 2932
rect 34428 2932 34512 2952
rect 34428 2924 34448 2932
rect 34456 2924 34484 2932
rect 34492 2924 34512 2932
rect 34548 2932 34632 2952
rect 34548 2924 34568 2932
rect 34576 2924 34604 2932
rect 34612 2924 34632 2932
rect 34668 2932 34752 2952
rect 34668 2924 34688 2932
rect 34696 2924 34724 2932
rect 34732 2924 34752 2932
rect 34788 2932 34872 2952
rect 34788 2924 34808 2932
rect 34816 2924 34844 2932
rect 34852 2924 34872 2932
rect 34908 2932 34992 2952
rect 34908 2924 34928 2932
rect 34936 2924 34964 2932
rect 34972 2924 34992 2932
rect 35028 2932 35112 2952
rect 35028 2924 35048 2932
rect 35056 2924 35084 2932
rect 35092 2924 35112 2932
rect 35148 2932 35232 2952
rect 35148 2924 35168 2932
rect 35176 2924 35204 2932
rect 35212 2924 35232 2932
rect 35268 2932 35352 2952
rect 35268 2924 35288 2932
rect 35296 2924 35324 2932
rect 35332 2924 35352 2932
rect 35388 2932 35472 2952
rect 35388 2924 35408 2932
rect 35416 2924 35444 2932
rect 35452 2924 35472 2932
rect 35508 2932 35592 2952
rect 35508 2924 35528 2932
rect 35536 2924 35564 2932
rect 35572 2924 35592 2932
rect 35628 2932 35712 2952
rect 35628 2924 35648 2932
rect 35656 2924 35684 2932
rect 35692 2924 35712 2932
rect 35748 2932 35832 2952
rect 35748 2924 35768 2932
rect 35776 2924 35804 2932
rect 35812 2924 35832 2932
rect 35868 2932 35952 2952
rect 35868 2924 35888 2932
rect 35896 2924 35924 2932
rect 35932 2924 35952 2932
rect 35988 2932 36072 2952
rect 35988 2924 36008 2932
rect 36016 2924 36044 2932
rect 36052 2924 36072 2932
rect 36108 2932 36192 2952
rect 36108 2924 36128 2932
rect 36136 2924 36164 2932
rect 36172 2924 36192 2932
rect 36228 2932 36312 2952
rect 36228 2924 36248 2932
rect 36256 2924 36284 2932
rect 36292 2924 36312 2932
rect 36348 2932 36432 2952
rect 36348 2924 36368 2932
rect 36376 2924 36404 2932
rect 36412 2924 36432 2932
rect 36468 2932 36552 2952
rect 36468 2924 36488 2932
rect 36496 2924 36524 2932
rect 36532 2924 36552 2932
rect 36588 2932 36672 2952
rect 36588 2924 36608 2932
rect 36616 2924 36644 2932
rect 36652 2924 36672 2932
rect 36708 2932 36792 2952
rect 36708 2924 36728 2932
rect 36736 2924 36764 2932
rect 36772 2924 36792 2932
rect 36828 2932 36912 2952
rect 36828 2924 36848 2932
rect 36856 2924 36884 2932
rect 36892 2924 36912 2932
rect 36948 2932 37032 2952
rect 36948 2924 36968 2932
rect 36976 2924 37004 2932
rect 37012 2924 37032 2932
rect 37068 2932 37152 2952
rect 37068 2924 37088 2932
rect 37096 2924 37124 2932
rect 37132 2924 37152 2932
rect 37188 2932 37272 2952
rect 37188 2924 37208 2932
rect 37216 2924 37244 2932
rect 37252 2924 37272 2932
rect 37308 2932 37392 2952
rect 37308 2924 37328 2932
rect 37336 2924 37364 2932
rect 37372 2924 37392 2932
rect 37428 2932 37512 2952
rect 37428 2924 37448 2932
rect 37456 2924 37484 2932
rect 37492 2924 37512 2932
rect 37548 2932 37632 2952
rect 37548 2924 37568 2932
rect 37576 2924 37604 2932
rect 37612 2924 37632 2932
rect 37668 2932 37752 2952
rect 37668 2924 37688 2932
rect 37696 2924 37724 2932
rect 37732 2924 37752 2932
rect 37788 2932 37872 2952
rect 37788 2924 37808 2932
rect 37816 2924 37844 2932
rect 37852 2924 37872 2932
rect 37908 2932 37992 2952
rect 37908 2924 37928 2932
rect 37936 2924 37964 2932
rect 37972 2924 37992 2932
rect 38028 2932 38112 2952
rect 38028 2924 38048 2932
rect 38056 2924 38084 2932
rect 38092 2924 38112 2932
rect 38148 2932 38232 2952
rect 38148 2924 38168 2932
rect 38176 2924 38204 2932
rect 38212 2924 38232 2932
rect 38268 2932 38352 2952
rect 38268 2924 38288 2932
rect 38296 2924 38324 2932
rect 38332 2924 38352 2932
rect 38388 2932 38472 2952
rect 38388 2924 38408 2932
rect 38416 2924 38444 2932
rect 38452 2924 38472 2932
rect 38508 2932 38592 2952
rect 38508 2924 38528 2932
rect 38536 2924 38564 2932
rect 38572 2924 38592 2932
rect 38628 2932 38712 2952
rect 38628 2924 38648 2932
rect 38656 2924 38684 2932
rect 38692 2924 38712 2932
rect 38748 2932 38832 2952
rect 38748 2924 38768 2932
rect 38776 2924 38804 2932
rect 38812 2924 38832 2932
rect 38868 2932 38952 2952
rect 38868 2924 38888 2932
rect 38896 2924 38924 2932
rect 38932 2924 38952 2932
rect 38988 2932 39072 2952
rect 38988 2924 39008 2932
rect 39016 2924 39044 2932
rect 39052 2924 39072 2932
rect 39108 2932 39192 2952
rect 39108 2924 39128 2932
rect 39136 2924 39164 2932
rect 39172 2924 39192 2932
rect 39228 2932 39312 2952
rect 39228 2924 39248 2932
rect 39256 2924 39284 2932
rect 39292 2924 39312 2932
rect 39348 2932 39432 2952
rect 39348 2924 39368 2932
rect 39376 2924 39404 2932
rect 39412 2924 39432 2932
rect 39468 2932 39552 2952
rect 39468 2924 39488 2932
rect 39496 2924 39524 2932
rect 39532 2924 39552 2932
rect 39588 2932 39672 2952
rect 39588 2924 39608 2932
rect 39616 2924 39644 2932
rect 39652 2924 39672 2932
rect 39708 2932 39792 2952
rect 39708 2924 39728 2932
rect 39736 2924 39764 2932
rect 39772 2924 39792 2932
rect 39828 2932 39912 2952
rect 39828 2924 39848 2932
rect 39856 2924 39884 2932
rect 39892 2924 39912 2932
rect 39948 2932 40032 2952
rect 39948 2924 39968 2932
rect 39976 2924 40004 2932
rect 40012 2924 40032 2932
rect 40068 2932 40152 2952
rect 40068 2924 40088 2932
rect 40096 2924 40124 2932
rect 40132 2924 40152 2932
rect 40188 2932 40272 2952
rect 40188 2924 40208 2932
rect 40216 2924 40244 2932
rect 40252 2924 40272 2932
rect 40308 2932 40392 2952
rect 40308 2924 40328 2932
rect 40336 2924 40364 2932
rect 40372 2924 40392 2932
rect 40428 2932 40512 2952
rect 40428 2924 40448 2932
rect 40456 2924 40484 2932
rect 40492 2924 40512 2932
rect 40548 2932 40632 2952
rect 40548 2924 40568 2932
rect 40576 2924 40604 2932
rect 40612 2924 40632 2932
rect 40668 2932 40752 2952
rect 40668 2924 40688 2932
rect 40696 2924 40724 2932
rect 40732 2924 40752 2932
rect 40788 2932 40872 2952
rect 40788 2924 40808 2932
rect 40816 2924 40844 2932
rect 40852 2924 40872 2932
rect 40908 2932 40992 2952
rect 40908 2924 40928 2932
rect 40936 2924 40964 2932
rect 40972 2924 40992 2932
rect 41028 2932 41112 2952
rect 41028 2924 41048 2932
rect 41056 2924 41084 2932
rect 41092 2924 41112 2932
rect 41148 2932 41232 2952
rect 41148 2924 41168 2932
rect 41176 2924 41204 2932
rect 41212 2924 41232 2932
rect 41268 2932 41352 2952
rect 41268 2924 41288 2932
rect 41296 2924 41324 2932
rect 41332 2924 41352 2932
rect 41388 2932 41472 2952
rect 41388 2924 41408 2932
rect 41416 2924 41444 2932
rect 41452 2924 41472 2932
rect 41508 2932 41592 2952
rect 41508 2924 41528 2932
rect 41536 2924 41564 2932
rect 41572 2924 41592 2932
rect 41628 2932 41712 2952
rect 41628 2924 41648 2932
rect 41656 2924 41684 2932
rect 41692 2924 41712 2932
rect 41748 2932 41832 2952
rect 41748 2924 41768 2932
rect 41776 2924 41804 2932
rect 41812 2924 41832 2932
rect 41868 2932 41952 2952
rect 41868 2924 41888 2932
rect 41896 2924 41924 2932
rect 41932 2924 41952 2932
rect 41988 2932 42072 2952
rect 41988 2924 42008 2932
rect 42016 2924 42044 2932
rect 42052 2924 42072 2932
rect 42108 2932 42192 2952
rect 42108 2924 42128 2932
rect 42136 2924 42164 2932
rect 42172 2924 42192 2932
rect 42228 2932 42312 2952
rect 42228 2924 42248 2932
rect 42256 2924 42284 2932
rect 42292 2924 42312 2932
rect 42348 2932 42432 2952
rect 42348 2924 42368 2932
rect 42376 2924 42404 2932
rect 42412 2924 42432 2932
rect 42468 2932 42552 2952
rect 42468 2924 42488 2932
rect 42496 2924 42524 2932
rect 42532 2924 42552 2932
rect 42588 2932 42672 2952
rect 42588 2924 42608 2932
rect 42616 2924 42644 2932
rect 42652 2924 42672 2932
rect 42708 2932 42792 2952
rect 42708 2924 42728 2932
rect 42736 2924 42764 2932
rect 42772 2924 42792 2932
rect 42828 2932 42912 2952
rect 42828 2924 42848 2932
rect 42856 2924 42884 2932
rect 42892 2924 42912 2932
rect 42948 2932 43032 2952
rect 42948 2924 42968 2932
rect 42976 2924 43004 2932
rect 43012 2924 43032 2932
rect 43068 2932 43152 2952
rect 43068 2924 43088 2932
rect 43096 2924 43124 2932
rect 43132 2924 43152 2932
rect 43188 2932 43272 2952
rect 43188 2924 43208 2932
rect 43216 2924 43244 2932
rect 43252 2924 43272 2932
rect 43308 2932 43392 2952
rect 43308 2924 43328 2932
rect 43336 2924 43364 2932
rect 43372 2924 43392 2932
rect 43428 2932 43512 2952
rect 43428 2924 43448 2932
rect 43456 2924 43484 2932
rect 43492 2924 43512 2932
rect 43548 2932 43632 2952
rect 43548 2924 43568 2932
rect 43576 2924 43604 2932
rect 43612 2924 43632 2932
rect 43668 2932 43752 2952
rect 43668 2924 43688 2932
rect 43696 2924 43724 2932
rect 43732 2924 43752 2932
rect 43788 2932 43872 2952
rect 43788 2924 43808 2932
rect 43816 2924 43844 2932
rect 43852 2924 43872 2932
rect 43908 2932 43992 2952
rect 43908 2924 43928 2932
rect 43936 2924 43964 2932
rect 43972 2924 43992 2932
rect 44028 2932 44112 2952
rect 44028 2924 44048 2932
rect 44056 2924 44084 2932
rect 44092 2924 44112 2932
rect 44148 2932 44232 2952
rect 44148 2924 44168 2932
rect 44176 2924 44204 2932
rect 44212 2924 44232 2932
rect 44268 2932 44352 2952
rect 44268 2924 44288 2932
rect 44296 2924 44324 2932
rect 44332 2924 44352 2932
rect 44388 2932 44472 2952
rect 44388 2924 44408 2932
rect 44416 2924 44444 2932
rect 44452 2924 44472 2932
rect 44508 2932 44592 2952
rect 44508 2924 44528 2932
rect 44536 2924 44564 2932
rect 44572 2924 44592 2932
rect 44628 2932 44712 2952
rect 44628 2924 44648 2932
rect 44656 2924 44684 2932
rect 44692 2924 44712 2932
rect 44748 2932 44832 2952
rect 44748 2924 44768 2932
rect 44776 2924 44804 2932
rect 44812 2924 44832 2932
rect 44868 2932 44952 2952
rect 44868 2924 44888 2932
rect 44896 2924 44924 2932
rect 44932 2924 44952 2932
rect 44988 2932 45072 2952
rect 44988 2924 45008 2932
rect 45016 2924 45044 2932
rect 45052 2924 45072 2932
rect 45108 2932 45192 2952
rect 45108 2924 45128 2932
rect 45136 2924 45164 2932
rect 45172 2924 45192 2932
rect 45228 2932 45312 2952
rect 45228 2924 45248 2932
rect 45256 2924 45284 2932
rect 45292 2924 45312 2932
rect 45348 2932 45432 2952
rect 45348 2924 45368 2932
rect 45376 2924 45404 2932
rect 45412 2924 45432 2932
rect 45468 2932 45552 2952
rect 45468 2924 45488 2932
rect 45496 2924 45524 2932
rect 45532 2924 45552 2932
rect 45588 2932 45672 2952
rect 45588 2924 45608 2932
rect 45616 2924 45644 2932
rect 45652 2924 45672 2932
rect 25936 2896 25992 2924
rect 26056 2896 26112 2924
rect 26176 2896 26232 2924
rect 26296 2896 26352 2924
rect 26416 2896 26472 2924
rect 26536 2896 26592 2924
rect 26656 2896 26712 2924
rect 26776 2896 26832 2924
rect 26896 2896 26952 2924
rect 27016 2896 27072 2924
rect 27136 2896 27192 2924
rect 27256 2896 27312 2924
rect 27376 2896 27432 2924
rect 27496 2896 27552 2924
rect 27616 2896 27672 2924
rect 27736 2896 27792 2924
rect 27856 2896 27912 2924
rect 27976 2896 28032 2924
rect 28096 2896 28152 2924
rect 28216 2896 28272 2924
rect 28336 2896 28392 2924
rect 28456 2896 28512 2924
rect 28576 2896 28632 2924
rect 28696 2896 28752 2924
rect 28816 2896 28872 2924
rect 28936 2896 28992 2924
rect 29056 2896 29112 2924
rect 29176 2896 29232 2924
rect 29296 2896 29352 2924
rect 29416 2896 29472 2924
rect 29536 2896 29592 2924
rect 29656 2896 29712 2924
rect 29776 2896 29832 2924
rect 29896 2896 29952 2924
rect 30016 2896 30072 2924
rect 30136 2896 30192 2924
rect 30256 2896 30312 2924
rect 30376 2896 30432 2924
rect 30496 2896 30552 2924
rect 30616 2896 30672 2924
rect 30736 2896 30792 2924
rect 30856 2896 30912 2924
rect 30976 2896 31032 2924
rect 31096 2896 31152 2924
rect 31216 2896 31272 2924
rect 31336 2896 31392 2924
rect 31456 2896 31512 2924
rect 31576 2896 31632 2924
rect 31696 2896 31752 2924
rect 31816 2896 31872 2924
rect 31936 2896 31992 2924
rect 32056 2896 32112 2924
rect 32176 2896 32232 2924
rect 32296 2896 32352 2924
rect 32416 2896 32472 2924
rect 32536 2896 32592 2924
rect 32656 2896 32712 2924
rect 32776 2896 32832 2924
rect 32896 2896 32952 2924
rect 33016 2896 33072 2924
rect 33136 2896 33192 2924
rect 33256 2896 33312 2924
rect 33376 2896 33432 2924
rect 33496 2896 33552 2924
rect 33616 2896 33672 2924
rect 33736 2896 33792 2924
rect 33856 2896 33912 2924
rect 33976 2896 34032 2924
rect 34096 2896 34152 2924
rect 34216 2896 34272 2924
rect 34336 2896 34392 2924
rect 34456 2896 34512 2924
rect 34576 2896 34632 2924
rect 34696 2896 34752 2924
rect 34816 2896 34872 2924
rect 34936 2896 34992 2924
rect 35056 2896 35112 2924
rect 35176 2896 35232 2924
rect 35296 2896 35352 2924
rect 35416 2896 35472 2924
rect 35536 2896 35592 2924
rect 35656 2896 35712 2924
rect 35776 2896 35832 2924
rect 35896 2896 35952 2924
rect 36016 2896 36072 2924
rect 36136 2896 36192 2924
rect 36256 2896 36312 2924
rect 36376 2896 36432 2924
rect 36496 2896 36552 2924
rect 36616 2896 36672 2924
rect 36736 2896 36792 2924
rect 36856 2896 36912 2924
rect 36976 2896 37032 2924
rect 37096 2896 37152 2924
rect 37216 2896 37272 2924
rect 37336 2896 37392 2924
rect 37456 2896 37512 2924
rect 37576 2896 37632 2924
rect 37696 2896 37752 2924
rect 37816 2896 37872 2924
rect 37936 2896 37992 2924
rect 38056 2896 38112 2924
rect 38176 2896 38232 2924
rect 38296 2896 38352 2924
rect 38416 2896 38472 2924
rect 38536 2896 38592 2924
rect 38656 2896 38712 2924
rect 38776 2896 38832 2924
rect 38896 2896 38952 2924
rect 39016 2896 39072 2924
rect 39136 2896 39192 2924
rect 39256 2896 39312 2924
rect 39376 2896 39432 2924
rect 39496 2896 39552 2924
rect 39616 2896 39672 2924
rect 39736 2896 39792 2924
rect 39856 2896 39912 2924
rect 39976 2896 40032 2924
rect 40096 2896 40152 2924
rect 40216 2896 40272 2924
rect 40336 2896 40392 2924
rect 40456 2896 40512 2924
rect 40576 2896 40632 2924
rect 40696 2896 40752 2924
rect 40816 2896 40872 2924
rect 40936 2896 40992 2924
rect 41056 2896 41112 2924
rect 41176 2896 41232 2924
rect 41296 2896 41352 2924
rect 41416 2896 41472 2924
rect 41536 2896 41592 2924
rect 41656 2896 41712 2924
rect 41776 2896 41832 2924
rect 41896 2896 41952 2924
rect 42016 2896 42072 2924
rect 42136 2896 42192 2924
rect 42256 2896 42312 2924
rect 42376 2896 42432 2924
rect 42496 2896 42552 2924
rect 42616 2896 42672 2924
rect 42736 2896 42792 2924
rect 42856 2896 42912 2924
rect 42976 2896 43032 2924
rect 43096 2896 43152 2924
rect 43216 2896 43272 2924
rect 43336 2896 43392 2924
rect 43456 2896 43512 2924
rect 43576 2896 43632 2924
rect 43696 2896 43752 2924
rect 43816 2896 43872 2924
rect 43936 2896 43992 2924
rect 44056 2896 44112 2924
rect 44176 2896 44232 2924
rect 44296 2896 44352 2924
rect 44416 2896 44472 2924
rect 44536 2896 44592 2924
rect 44656 2896 44712 2924
rect 44776 2896 44832 2924
rect 44896 2896 44952 2924
rect 45016 2896 45072 2924
rect 45136 2896 45192 2924
rect 45256 2896 45312 2924
rect 45376 2896 45432 2924
rect 45496 2896 45552 2924
rect 45616 2896 45672 2924
rect 25908 2752 25992 2772
rect 25908 2744 25928 2752
rect 25936 2744 25964 2752
rect 25972 2744 25992 2752
rect 26028 2752 26112 2772
rect 26028 2744 26048 2752
rect 26056 2744 26084 2752
rect 26092 2744 26112 2752
rect 26148 2752 26232 2772
rect 26148 2744 26168 2752
rect 26176 2744 26204 2752
rect 26212 2744 26232 2752
rect 26268 2752 26352 2772
rect 26268 2744 26288 2752
rect 26296 2744 26324 2752
rect 26332 2744 26352 2752
rect 26388 2752 26472 2772
rect 26388 2744 26408 2752
rect 26416 2744 26444 2752
rect 26452 2744 26472 2752
rect 26508 2752 26592 2772
rect 26508 2744 26528 2752
rect 26536 2744 26564 2752
rect 26572 2744 26592 2752
rect 26628 2752 26712 2772
rect 26628 2744 26648 2752
rect 26656 2744 26684 2752
rect 26692 2744 26712 2752
rect 26748 2752 26832 2772
rect 26748 2744 26768 2752
rect 26776 2744 26804 2752
rect 26812 2744 26832 2752
rect 26868 2752 26952 2772
rect 26868 2744 26888 2752
rect 26896 2744 26924 2752
rect 26932 2744 26952 2752
rect 26988 2752 27072 2772
rect 26988 2744 27008 2752
rect 27016 2744 27044 2752
rect 27052 2744 27072 2752
rect 27108 2752 27192 2772
rect 27108 2744 27128 2752
rect 27136 2744 27164 2752
rect 27172 2744 27192 2752
rect 27228 2752 27312 2772
rect 27228 2744 27248 2752
rect 27256 2744 27284 2752
rect 27292 2744 27312 2752
rect 27348 2752 27432 2772
rect 27348 2744 27368 2752
rect 27376 2744 27404 2752
rect 27412 2744 27432 2752
rect 27468 2752 27552 2772
rect 27468 2744 27488 2752
rect 27496 2744 27524 2752
rect 27532 2744 27552 2752
rect 27588 2752 27672 2772
rect 27588 2744 27608 2752
rect 27616 2744 27644 2752
rect 27652 2744 27672 2752
rect 27708 2752 27792 2772
rect 27708 2744 27728 2752
rect 27736 2744 27764 2752
rect 27772 2744 27792 2752
rect 27828 2752 27912 2772
rect 27828 2744 27848 2752
rect 27856 2744 27884 2752
rect 27892 2744 27912 2752
rect 27948 2752 28032 2772
rect 27948 2744 27968 2752
rect 27976 2744 28004 2752
rect 28012 2744 28032 2752
rect 28068 2752 28152 2772
rect 28068 2744 28088 2752
rect 28096 2744 28124 2752
rect 28132 2744 28152 2752
rect 28188 2752 28272 2772
rect 28188 2744 28208 2752
rect 28216 2744 28244 2752
rect 28252 2744 28272 2752
rect 28308 2752 28392 2772
rect 28308 2744 28328 2752
rect 28336 2744 28364 2752
rect 28372 2744 28392 2752
rect 28428 2752 28512 2772
rect 28428 2744 28448 2752
rect 28456 2744 28484 2752
rect 28492 2744 28512 2752
rect 28548 2752 28632 2772
rect 28548 2744 28568 2752
rect 28576 2744 28604 2752
rect 28612 2744 28632 2752
rect 28668 2752 28752 2772
rect 28668 2744 28688 2752
rect 28696 2744 28724 2752
rect 28732 2744 28752 2752
rect 28788 2752 28872 2772
rect 28788 2744 28808 2752
rect 28816 2744 28844 2752
rect 28852 2744 28872 2752
rect 28908 2752 28992 2772
rect 28908 2744 28928 2752
rect 28936 2744 28964 2752
rect 28972 2744 28992 2752
rect 29028 2752 29112 2772
rect 29028 2744 29048 2752
rect 29056 2744 29084 2752
rect 29092 2744 29112 2752
rect 29148 2752 29232 2772
rect 29148 2744 29168 2752
rect 29176 2744 29204 2752
rect 29212 2744 29232 2752
rect 29268 2752 29352 2772
rect 29268 2744 29288 2752
rect 29296 2744 29324 2752
rect 29332 2744 29352 2752
rect 29388 2752 29472 2772
rect 29388 2744 29408 2752
rect 29416 2744 29444 2752
rect 29452 2744 29472 2752
rect 29508 2752 29592 2772
rect 29508 2744 29528 2752
rect 29536 2744 29564 2752
rect 29572 2744 29592 2752
rect 29628 2752 29712 2772
rect 29628 2744 29648 2752
rect 29656 2744 29684 2752
rect 29692 2744 29712 2752
rect 29748 2752 29832 2772
rect 29748 2744 29768 2752
rect 29776 2744 29804 2752
rect 29812 2744 29832 2752
rect 29868 2752 29952 2772
rect 29868 2744 29888 2752
rect 29896 2744 29924 2752
rect 29932 2744 29952 2752
rect 29988 2752 30072 2772
rect 29988 2744 30008 2752
rect 30016 2744 30044 2752
rect 30052 2744 30072 2752
rect 30108 2752 30192 2772
rect 30108 2744 30128 2752
rect 30136 2744 30164 2752
rect 30172 2744 30192 2752
rect 30228 2752 30312 2772
rect 30228 2744 30248 2752
rect 30256 2744 30284 2752
rect 30292 2744 30312 2752
rect 30348 2752 30432 2772
rect 30348 2744 30368 2752
rect 30376 2744 30404 2752
rect 30412 2744 30432 2752
rect 30468 2752 30552 2772
rect 30468 2744 30488 2752
rect 30496 2744 30524 2752
rect 30532 2744 30552 2752
rect 30588 2752 30672 2772
rect 30588 2744 30608 2752
rect 30616 2744 30644 2752
rect 30652 2744 30672 2752
rect 30708 2752 30792 2772
rect 30708 2744 30728 2752
rect 30736 2744 30764 2752
rect 30772 2744 30792 2752
rect 30828 2752 30912 2772
rect 30828 2744 30848 2752
rect 30856 2744 30884 2752
rect 30892 2744 30912 2752
rect 30948 2752 31032 2772
rect 30948 2744 30968 2752
rect 30976 2744 31004 2752
rect 31012 2744 31032 2752
rect 31068 2752 31152 2772
rect 31068 2744 31088 2752
rect 31096 2744 31124 2752
rect 31132 2744 31152 2752
rect 31188 2752 31272 2772
rect 31188 2744 31208 2752
rect 31216 2744 31244 2752
rect 31252 2744 31272 2752
rect 31308 2752 31392 2772
rect 31308 2744 31328 2752
rect 31336 2744 31364 2752
rect 31372 2744 31392 2752
rect 31428 2752 31512 2772
rect 31428 2744 31448 2752
rect 31456 2744 31484 2752
rect 31492 2744 31512 2752
rect 31548 2752 31632 2772
rect 31548 2744 31568 2752
rect 31576 2744 31604 2752
rect 31612 2744 31632 2752
rect 31668 2752 31752 2772
rect 31668 2744 31688 2752
rect 31696 2744 31724 2752
rect 31732 2744 31752 2752
rect 31788 2752 31872 2772
rect 31788 2744 31808 2752
rect 31816 2744 31844 2752
rect 31852 2744 31872 2752
rect 31908 2752 31992 2772
rect 31908 2744 31928 2752
rect 31936 2744 31964 2752
rect 31972 2744 31992 2752
rect 32028 2752 32112 2772
rect 32028 2744 32048 2752
rect 32056 2744 32084 2752
rect 32092 2744 32112 2752
rect 32148 2752 32232 2772
rect 32148 2744 32168 2752
rect 32176 2744 32204 2752
rect 32212 2744 32232 2752
rect 32268 2752 32352 2772
rect 32268 2744 32288 2752
rect 32296 2744 32324 2752
rect 32332 2744 32352 2752
rect 32388 2752 32472 2772
rect 32388 2744 32408 2752
rect 32416 2744 32444 2752
rect 32452 2744 32472 2752
rect 32508 2752 32592 2772
rect 32508 2744 32528 2752
rect 32536 2744 32564 2752
rect 32572 2744 32592 2752
rect 32628 2752 32712 2772
rect 32628 2744 32648 2752
rect 32656 2744 32684 2752
rect 32692 2744 32712 2752
rect 32748 2752 32832 2772
rect 32748 2744 32768 2752
rect 32776 2744 32804 2752
rect 32812 2744 32832 2752
rect 32868 2752 32952 2772
rect 32868 2744 32888 2752
rect 32896 2744 32924 2752
rect 32932 2744 32952 2752
rect 32988 2752 33072 2772
rect 32988 2744 33008 2752
rect 33016 2744 33044 2752
rect 33052 2744 33072 2752
rect 33108 2752 33192 2772
rect 33108 2744 33128 2752
rect 33136 2744 33164 2752
rect 33172 2744 33192 2752
rect 33228 2752 33312 2772
rect 33228 2744 33248 2752
rect 33256 2744 33284 2752
rect 33292 2744 33312 2752
rect 33348 2752 33432 2772
rect 33348 2744 33368 2752
rect 33376 2744 33404 2752
rect 33412 2744 33432 2752
rect 33468 2752 33552 2772
rect 33468 2744 33488 2752
rect 33496 2744 33524 2752
rect 33532 2744 33552 2752
rect 33588 2752 33672 2772
rect 33588 2744 33608 2752
rect 33616 2744 33644 2752
rect 33652 2744 33672 2752
rect 33708 2752 33792 2772
rect 33708 2744 33728 2752
rect 33736 2744 33764 2752
rect 33772 2744 33792 2752
rect 33828 2752 33912 2772
rect 33828 2744 33848 2752
rect 33856 2744 33884 2752
rect 33892 2744 33912 2752
rect 33948 2752 34032 2772
rect 33948 2744 33968 2752
rect 33976 2744 34004 2752
rect 34012 2744 34032 2752
rect 34068 2752 34152 2772
rect 34068 2744 34088 2752
rect 34096 2744 34124 2752
rect 34132 2744 34152 2752
rect 34188 2752 34272 2772
rect 34188 2744 34208 2752
rect 34216 2744 34244 2752
rect 34252 2744 34272 2752
rect 34308 2752 34392 2772
rect 34308 2744 34328 2752
rect 34336 2744 34364 2752
rect 34372 2744 34392 2752
rect 34428 2752 34512 2772
rect 34428 2744 34448 2752
rect 34456 2744 34484 2752
rect 34492 2744 34512 2752
rect 34548 2752 34632 2772
rect 34548 2744 34568 2752
rect 34576 2744 34604 2752
rect 34612 2744 34632 2752
rect 34668 2752 34752 2772
rect 34668 2744 34688 2752
rect 34696 2744 34724 2752
rect 34732 2744 34752 2752
rect 34788 2752 34872 2772
rect 34788 2744 34808 2752
rect 34816 2744 34844 2752
rect 34852 2744 34872 2752
rect 34908 2752 34992 2772
rect 34908 2744 34928 2752
rect 34936 2744 34964 2752
rect 34972 2744 34992 2752
rect 35028 2752 35112 2772
rect 35028 2744 35048 2752
rect 35056 2744 35084 2752
rect 35092 2744 35112 2752
rect 35148 2752 35232 2772
rect 35148 2744 35168 2752
rect 35176 2744 35204 2752
rect 35212 2744 35232 2752
rect 35268 2752 35352 2772
rect 35268 2744 35288 2752
rect 35296 2744 35324 2752
rect 35332 2744 35352 2752
rect 35388 2752 35472 2772
rect 35388 2744 35408 2752
rect 35416 2744 35444 2752
rect 35452 2744 35472 2752
rect 35508 2752 35592 2772
rect 35508 2744 35528 2752
rect 35536 2744 35564 2752
rect 35572 2744 35592 2752
rect 35628 2752 35712 2772
rect 35628 2744 35648 2752
rect 35656 2744 35684 2752
rect 35692 2744 35712 2752
rect 35748 2752 35832 2772
rect 35748 2744 35768 2752
rect 35776 2744 35804 2752
rect 35812 2744 35832 2752
rect 35868 2752 35952 2772
rect 35868 2744 35888 2752
rect 35896 2744 35924 2752
rect 35932 2744 35952 2752
rect 35988 2752 36072 2772
rect 35988 2744 36008 2752
rect 36016 2744 36044 2752
rect 36052 2744 36072 2752
rect 36108 2752 36192 2772
rect 36108 2744 36128 2752
rect 36136 2744 36164 2752
rect 36172 2744 36192 2752
rect 36228 2752 36312 2772
rect 36228 2744 36248 2752
rect 36256 2744 36284 2752
rect 36292 2744 36312 2752
rect 36348 2752 36432 2772
rect 36348 2744 36368 2752
rect 36376 2744 36404 2752
rect 36412 2744 36432 2752
rect 36468 2752 36552 2772
rect 36468 2744 36488 2752
rect 36496 2744 36524 2752
rect 36532 2744 36552 2752
rect 36588 2752 36672 2772
rect 36588 2744 36608 2752
rect 36616 2744 36644 2752
rect 36652 2744 36672 2752
rect 36708 2752 36792 2772
rect 36708 2744 36728 2752
rect 36736 2744 36764 2752
rect 36772 2744 36792 2752
rect 36828 2752 36912 2772
rect 36828 2744 36848 2752
rect 36856 2744 36884 2752
rect 36892 2744 36912 2752
rect 36948 2752 37032 2772
rect 36948 2744 36968 2752
rect 36976 2744 37004 2752
rect 37012 2744 37032 2752
rect 37068 2752 37152 2772
rect 37068 2744 37088 2752
rect 37096 2744 37124 2752
rect 37132 2744 37152 2752
rect 37188 2752 37272 2772
rect 37188 2744 37208 2752
rect 37216 2744 37244 2752
rect 37252 2744 37272 2752
rect 37308 2752 37392 2772
rect 37308 2744 37328 2752
rect 37336 2744 37364 2752
rect 37372 2744 37392 2752
rect 37428 2752 37512 2772
rect 37428 2744 37448 2752
rect 37456 2744 37484 2752
rect 37492 2744 37512 2752
rect 37548 2752 37632 2772
rect 37548 2744 37568 2752
rect 37576 2744 37604 2752
rect 37612 2744 37632 2752
rect 37668 2752 37752 2772
rect 37668 2744 37688 2752
rect 37696 2744 37724 2752
rect 37732 2744 37752 2752
rect 37788 2752 37872 2772
rect 37788 2744 37808 2752
rect 37816 2744 37844 2752
rect 37852 2744 37872 2752
rect 37908 2752 37992 2772
rect 37908 2744 37928 2752
rect 37936 2744 37964 2752
rect 37972 2744 37992 2752
rect 38028 2752 38112 2772
rect 38028 2744 38048 2752
rect 38056 2744 38084 2752
rect 38092 2744 38112 2752
rect 38148 2752 38232 2772
rect 38148 2744 38168 2752
rect 38176 2744 38204 2752
rect 38212 2744 38232 2752
rect 38268 2752 38352 2772
rect 38268 2744 38288 2752
rect 38296 2744 38324 2752
rect 38332 2744 38352 2752
rect 38388 2752 38472 2772
rect 38388 2744 38408 2752
rect 38416 2744 38444 2752
rect 38452 2744 38472 2752
rect 38508 2752 38592 2772
rect 38508 2744 38528 2752
rect 38536 2744 38564 2752
rect 38572 2744 38592 2752
rect 38628 2752 38712 2772
rect 38628 2744 38648 2752
rect 38656 2744 38684 2752
rect 38692 2744 38712 2752
rect 38748 2752 38832 2772
rect 38748 2744 38768 2752
rect 38776 2744 38804 2752
rect 38812 2744 38832 2752
rect 38868 2752 38952 2772
rect 38868 2744 38888 2752
rect 38896 2744 38924 2752
rect 38932 2744 38952 2752
rect 38988 2752 39072 2772
rect 38988 2744 39008 2752
rect 39016 2744 39044 2752
rect 39052 2744 39072 2752
rect 39108 2752 39192 2772
rect 39108 2744 39128 2752
rect 39136 2744 39164 2752
rect 39172 2744 39192 2752
rect 39228 2752 39312 2772
rect 39228 2744 39248 2752
rect 39256 2744 39284 2752
rect 39292 2744 39312 2752
rect 39348 2752 39432 2772
rect 39348 2744 39368 2752
rect 39376 2744 39404 2752
rect 39412 2744 39432 2752
rect 39468 2752 39552 2772
rect 39468 2744 39488 2752
rect 39496 2744 39524 2752
rect 39532 2744 39552 2752
rect 39588 2752 39672 2772
rect 39588 2744 39608 2752
rect 39616 2744 39644 2752
rect 39652 2744 39672 2752
rect 39708 2752 39792 2772
rect 39708 2744 39728 2752
rect 39736 2744 39764 2752
rect 39772 2744 39792 2752
rect 39828 2752 39912 2772
rect 39828 2744 39848 2752
rect 39856 2744 39884 2752
rect 39892 2744 39912 2752
rect 39948 2752 40032 2772
rect 39948 2744 39968 2752
rect 39976 2744 40004 2752
rect 40012 2744 40032 2752
rect 40068 2752 40152 2772
rect 40068 2744 40088 2752
rect 40096 2744 40124 2752
rect 40132 2744 40152 2752
rect 40188 2752 40272 2772
rect 40188 2744 40208 2752
rect 40216 2744 40244 2752
rect 40252 2744 40272 2752
rect 40308 2752 40392 2772
rect 40308 2744 40328 2752
rect 40336 2744 40364 2752
rect 40372 2744 40392 2752
rect 40428 2752 40512 2772
rect 40428 2744 40448 2752
rect 40456 2744 40484 2752
rect 40492 2744 40512 2752
rect 40548 2752 40632 2772
rect 40548 2744 40568 2752
rect 40576 2744 40604 2752
rect 40612 2744 40632 2752
rect 40668 2752 40752 2772
rect 40668 2744 40688 2752
rect 40696 2744 40724 2752
rect 40732 2744 40752 2752
rect 40788 2752 40872 2772
rect 40788 2744 40808 2752
rect 40816 2744 40844 2752
rect 40852 2744 40872 2752
rect 40908 2752 40992 2772
rect 40908 2744 40928 2752
rect 40936 2744 40964 2752
rect 40972 2744 40992 2752
rect 41028 2752 41112 2772
rect 41028 2744 41048 2752
rect 41056 2744 41084 2752
rect 41092 2744 41112 2752
rect 41148 2752 41232 2772
rect 41148 2744 41168 2752
rect 41176 2744 41204 2752
rect 41212 2744 41232 2752
rect 41268 2752 41352 2772
rect 41268 2744 41288 2752
rect 41296 2744 41324 2752
rect 41332 2744 41352 2752
rect 41388 2752 41472 2772
rect 41388 2744 41408 2752
rect 41416 2744 41444 2752
rect 41452 2744 41472 2752
rect 41508 2752 41592 2772
rect 41508 2744 41528 2752
rect 41536 2744 41564 2752
rect 41572 2744 41592 2752
rect 41628 2752 41712 2772
rect 41628 2744 41648 2752
rect 41656 2744 41684 2752
rect 41692 2744 41712 2752
rect 41748 2752 41832 2772
rect 41748 2744 41768 2752
rect 41776 2744 41804 2752
rect 41812 2744 41832 2752
rect 41868 2752 41952 2772
rect 41868 2744 41888 2752
rect 41896 2744 41924 2752
rect 41932 2744 41952 2752
rect 41988 2752 42072 2772
rect 41988 2744 42008 2752
rect 42016 2744 42044 2752
rect 42052 2744 42072 2752
rect 42108 2752 42192 2772
rect 42108 2744 42128 2752
rect 42136 2744 42164 2752
rect 42172 2744 42192 2752
rect 42228 2752 42312 2772
rect 42228 2744 42248 2752
rect 42256 2744 42284 2752
rect 42292 2744 42312 2752
rect 42348 2752 42432 2772
rect 42348 2744 42368 2752
rect 42376 2744 42404 2752
rect 42412 2744 42432 2752
rect 42468 2752 42552 2772
rect 42468 2744 42488 2752
rect 42496 2744 42524 2752
rect 42532 2744 42552 2752
rect 42588 2752 42672 2772
rect 42588 2744 42608 2752
rect 42616 2744 42644 2752
rect 42652 2744 42672 2752
rect 42708 2752 42792 2772
rect 42708 2744 42728 2752
rect 42736 2744 42764 2752
rect 42772 2744 42792 2752
rect 42828 2752 42912 2772
rect 42828 2744 42848 2752
rect 42856 2744 42884 2752
rect 42892 2744 42912 2752
rect 42948 2752 43032 2772
rect 42948 2744 42968 2752
rect 42976 2744 43004 2752
rect 43012 2744 43032 2752
rect 43068 2752 43152 2772
rect 43068 2744 43088 2752
rect 43096 2744 43124 2752
rect 43132 2744 43152 2752
rect 43188 2752 43272 2772
rect 43188 2744 43208 2752
rect 43216 2744 43244 2752
rect 43252 2744 43272 2752
rect 43308 2752 43392 2772
rect 43308 2744 43328 2752
rect 43336 2744 43364 2752
rect 43372 2744 43392 2752
rect 43428 2752 43512 2772
rect 43428 2744 43448 2752
rect 43456 2744 43484 2752
rect 43492 2744 43512 2752
rect 43548 2752 43632 2772
rect 43548 2744 43568 2752
rect 43576 2744 43604 2752
rect 43612 2744 43632 2752
rect 43668 2752 43752 2772
rect 43668 2744 43688 2752
rect 43696 2744 43724 2752
rect 43732 2744 43752 2752
rect 43788 2752 43872 2772
rect 43788 2744 43808 2752
rect 43816 2744 43844 2752
rect 43852 2744 43872 2752
rect 43908 2752 43992 2772
rect 43908 2744 43928 2752
rect 43936 2744 43964 2752
rect 43972 2744 43992 2752
rect 44028 2752 44112 2772
rect 44028 2744 44048 2752
rect 44056 2744 44084 2752
rect 44092 2744 44112 2752
rect 44148 2752 44232 2772
rect 44148 2744 44168 2752
rect 44176 2744 44204 2752
rect 44212 2744 44232 2752
rect 44268 2752 44352 2772
rect 44268 2744 44288 2752
rect 44296 2744 44324 2752
rect 44332 2744 44352 2752
rect 44388 2752 44472 2772
rect 44388 2744 44408 2752
rect 44416 2744 44444 2752
rect 44452 2744 44472 2752
rect 44508 2752 44592 2772
rect 44508 2744 44528 2752
rect 44536 2744 44564 2752
rect 44572 2744 44592 2752
rect 44628 2752 44712 2772
rect 44628 2744 44648 2752
rect 44656 2744 44684 2752
rect 44692 2744 44712 2752
rect 44748 2752 44832 2772
rect 44748 2744 44768 2752
rect 44776 2744 44804 2752
rect 44812 2744 44832 2752
rect 44868 2752 44952 2772
rect 44868 2744 44888 2752
rect 44896 2744 44924 2752
rect 44932 2744 44952 2752
rect 44988 2752 45072 2772
rect 44988 2744 45008 2752
rect 45016 2744 45044 2752
rect 45052 2744 45072 2752
rect 45108 2752 45192 2772
rect 45108 2744 45128 2752
rect 45136 2744 45164 2752
rect 45172 2744 45192 2752
rect 45228 2752 45312 2772
rect 45228 2744 45248 2752
rect 45256 2744 45284 2752
rect 45292 2744 45312 2752
rect 45348 2752 45432 2772
rect 45348 2744 45368 2752
rect 45376 2744 45404 2752
rect 45412 2744 45432 2752
rect 45468 2752 45552 2772
rect 45468 2744 45488 2752
rect 45496 2744 45524 2752
rect 45532 2744 45552 2752
rect 45588 2752 45672 2772
rect 45588 2744 45608 2752
rect 45616 2744 45644 2752
rect 45652 2744 45672 2752
rect 25936 2716 25992 2744
rect 26056 2716 26112 2744
rect 26176 2716 26232 2744
rect 26296 2716 26352 2744
rect 26416 2716 26472 2744
rect 26536 2716 26592 2744
rect 26656 2716 26712 2744
rect 26776 2716 26832 2744
rect 26896 2716 26952 2744
rect 27016 2716 27072 2744
rect 27136 2716 27192 2744
rect 27256 2716 27312 2744
rect 27376 2716 27432 2744
rect 27496 2716 27552 2744
rect 27616 2716 27672 2744
rect 27736 2716 27792 2744
rect 27856 2716 27912 2744
rect 27976 2716 28032 2744
rect 28096 2716 28152 2744
rect 28216 2716 28272 2744
rect 28336 2716 28392 2744
rect 28456 2716 28512 2744
rect 28576 2716 28632 2744
rect 28696 2716 28752 2744
rect 28816 2716 28872 2744
rect 28936 2716 28992 2744
rect 29056 2716 29112 2744
rect 29176 2716 29232 2744
rect 29296 2716 29352 2744
rect 29416 2716 29472 2744
rect 29536 2716 29592 2744
rect 29656 2716 29712 2744
rect 29776 2716 29832 2744
rect 29896 2716 29952 2744
rect 30016 2716 30072 2744
rect 30136 2716 30192 2744
rect 30256 2716 30312 2744
rect 30376 2716 30432 2744
rect 30496 2716 30552 2744
rect 30616 2716 30672 2744
rect 30736 2716 30792 2744
rect 30856 2716 30912 2744
rect 30976 2716 31032 2744
rect 31096 2716 31152 2744
rect 31216 2716 31272 2744
rect 31336 2716 31392 2744
rect 31456 2716 31512 2744
rect 31576 2716 31632 2744
rect 31696 2716 31752 2744
rect 31816 2716 31872 2744
rect 31936 2716 31992 2744
rect 32056 2716 32112 2744
rect 32176 2716 32232 2744
rect 32296 2716 32352 2744
rect 32416 2716 32472 2744
rect 32536 2716 32592 2744
rect 32656 2716 32712 2744
rect 32776 2716 32832 2744
rect 32896 2716 32952 2744
rect 33016 2716 33072 2744
rect 33136 2716 33192 2744
rect 33256 2716 33312 2744
rect 33376 2716 33432 2744
rect 33496 2716 33552 2744
rect 33616 2716 33672 2744
rect 33736 2716 33792 2744
rect 33856 2716 33912 2744
rect 33976 2716 34032 2744
rect 34096 2716 34152 2744
rect 34216 2716 34272 2744
rect 34336 2716 34392 2744
rect 34456 2716 34512 2744
rect 34576 2716 34632 2744
rect 34696 2716 34752 2744
rect 34816 2716 34872 2744
rect 34936 2716 34992 2744
rect 35056 2716 35112 2744
rect 35176 2716 35232 2744
rect 35296 2716 35352 2744
rect 35416 2716 35472 2744
rect 35536 2716 35592 2744
rect 35656 2716 35712 2744
rect 35776 2716 35832 2744
rect 35896 2716 35952 2744
rect 36016 2716 36072 2744
rect 36136 2716 36192 2744
rect 36256 2716 36312 2744
rect 36376 2716 36432 2744
rect 36496 2716 36552 2744
rect 36616 2716 36672 2744
rect 36736 2716 36792 2744
rect 36856 2716 36912 2744
rect 36976 2716 37032 2744
rect 37096 2716 37152 2744
rect 37216 2716 37272 2744
rect 37336 2716 37392 2744
rect 37456 2716 37512 2744
rect 37576 2716 37632 2744
rect 37696 2716 37752 2744
rect 37816 2716 37872 2744
rect 37936 2716 37992 2744
rect 38056 2716 38112 2744
rect 38176 2716 38232 2744
rect 38296 2716 38352 2744
rect 38416 2716 38472 2744
rect 38536 2716 38592 2744
rect 38656 2716 38712 2744
rect 38776 2716 38832 2744
rect 38896 2716 38952 2744
rect 39016 2716 39072 2744
rect 39136 2716 39192 2744
rect 39256 2716 39312 2744
rect 39376 2716 39432 2744
rect 39496 2716 39552 2744
rect 39616 2716 39672 2744
rect 39736 2716 39792 2744
rect 39856 2716 39912 2744
rect 39976 2716 40032 2744
rect 40096 2716 40152 2744
rect 40216 2716 40272 2744
rect 40336 2716 40392 2744
rect 40456 2716 40512 2744
rect 40576 2716 40632 2744
rect 40696 2716 40752 2744
rect 40816 2716 40872 2744
rect 40936 2716 40992 2744
rect 41056 2716 41112 2744
rect 41176 2716 41232 2744
rect 41296 2716 41352 2744
rect 41416 2716 41472 2744
rect 41536 2716 41592 2744
rect 41656 2716 41712 2744
rect 41776 2716 41832 2744
rect 41896 2716 41952 2744
rect 42016 2716 42072 2744
rect 42136 2716 42192 2744
rect 42256 2716 42312 2744
rect 42376 2716 42432 2744
rect 42496 2716 42552 2744
rect 42616 2716 42672 2744
rect 42736 2716 42792 2744
rect 42856 2716 42912 2744
rect 42976 2716 43032 2744
rect 43096 2716 43152 2744
rect 43216 2716 43272 2744
rect 43336 2716 43392 2744
rect 43456 2716 43512 2744
rect 43576 2716 43632 2744
rect 43696 2716 43752 2744
rect 43816 2716 43872 2744
rect 43936 2716 43992 2744
rect 44056 2716 44112 2744
rect 44176 2716 44232 2744
rect 44296 2716 44352 2744
rect 44416 2716 44472 2744
rect 44536 2716 44592 2744
rect 44656 2716 44712 2744
rect 44776 2716 44832 2744
rect 44896 2716 44952 2744
rect 45016 2716 45072 2744
rect 45136 2716 45192 2744
rect 45256 2716 45312 2744
rect 45376 2716 45432 2744
rect 45496 2716 45552 2744
rect 45616 2716 45672 2744
rect 25908 2572 25992 2592
rect 25908 2564 25928 2572
rect 25936 2564 25964 2572
rect 25972 2564 25992 2572
rect 26028 2572 26112 2592
rect 26028 2564 26048 2572
rect 26056 2564 26084 2572
rect 26092 2564 26112 2572
rect 26148 2572 26232 2592
rect 26148 2564 26168 2572
rect 26176 2564 26204 2572
rect 26212 2564 26232 2572
rect 26268 2572 26352 2592
rect 26268 2564 26288 2572
rect 26296 2564 26324 2572
rect 26332 2564 26352 2572
rect 26388 2572 26472 2592
rect 26388 2564 26408 2572
rect 26416 2564 26444 2572
rect 26452 2564 26472 2572
rect 26508 2572 26592 2592
rect 26508 2564 26528 2572
rect 26536 2564 26564 2572
rect 26572 2564 26592 2572
rect 26628 2572 26712 2592
rect 26628 2564 26648 2572
rect 26656 2564 26684 2572
rect 26692 2564 26712 2572
rect 26748 2572 26832 2592
rect 26748 2564 26768 2572
rect 26776 2564 26804 2572
rect 26812 2564 26832 2572
rect 26868 2572 26952 2592
rect 26868 2564 26888 2572
rect 26896 2564 26924 2572
rect 26932 2564 26952 2572
rect 26988 2572 27072 2592
rect 26988 2564 27008 2572
rect 27016 2564 27044 2572
rect 27052 2564 27072 2572
rect 27108 2572 27192 2592
rect 27108 2564 27128 2572
rect 27136 2564 27164 2572
rect 27172 2564 27192 2572
rect 27228 2572 27312 2592
rect 27228 2564 27248 2572
rect 27256 2564 27284 2572
rect 27292 2564 27312 2572
rect 27348 2572 27432 2592
rect 27348 2564 27368 2572
rect 27376 2564 27404 2572
rect 27412 2564 27432 2572
rect 27468 2572 27552 2592
rect 27468 2564 27488 2572
rect 27496 2564 27524 2572
rect 27532 2564 27552 2572
rect 27588 2572 27672 2592
rect 27588 2564 27608 2572
rect 27616 2564 27644 2572
rect 27652 2564 27672 2572
rect 27708 2572 27792 2592
rect 27708 2564 27728 2572
rect 27736 2564 27764 2572
rect 27772 2564 27792 2572
rect 27828 2572 27912 2592
rect 27828 2564 27848 2572
rect 27856 2564 27884 2572
rect 27892 2564 27912 2572
rect 27948 2572 28032 2592
rect 27948 2564 27968 2572
rect 27976 2564 28004 2572
rect 28012 2564 28032 2572
rect 28068 2572 28152 2592
rect 28068 2564 28088 2572
rect 28096 2564 28124 2572
rect 28132 2564 28152 2572
rect 28188 2572 28272 2592
rect 28188 2564 28208 2572
rect 28216 2564 28244 2572
rect 28252 2564 28272 2572
rect 28308 2572 28392 2592
rect 28308 2564 28328 2572
rect 28336 2564 28364 2572
rect 28372 2564 28392 2572
rect 28428 2572 28512 2592
rect 28428 2564 28448 2572
rect 28456 2564 28484 2572
rect 28492 2564 28512 2572
rect 28548 2572 28632 2592
rect 28548 2564 28568 2572
rect 28576 2564 28604 2572
rect 28612 2564 28632 2572
rect 28668 2572 28752 2592
rect 28668 2564 28688 2572
rect 28696 2564 28724 2572
rect 28732 2564 28752 2572
rect 28788 2572 28872 2592
rect 28788 2564 28808 2572
rect 28816 2564 28844 2572
rect 28852 2564 28872 2572
rect 28908 2572 28992 2592
rect 28908 2564 28928 2572
rect 28936 2564 28964 2572
rect 28972 2564 28992 2572
rect 29028 2572 29112 2592
rect 29028 2564 29048 2572
rect 29056 2564 29084 2572
rect 29092 2564 29112 2572
rect 29148 2572 29232 2592
rect 29148 2564 29168 2572
rect 29176 2564 29204 2572
rect 29212 2564 29232 2572
rect 29268 2572 29352 2592
rect 29268 2564 29288 2572
rect 29296 2564 29324 2572
rect 29332 2564 29352 2572
rect 29388 2572 29472 2592
rect 29388 2564 29408 2572
rect 29416 2564 29444 2572
rect 29452 2564 29472 2572
rect 29508 2572 29592 2592
rect 29508 2564 29528 2572
rect 29536 2564 29564 2572
rect 29572 2564 29592 2572
rect 29628 2572 29712 2592
rect 29628 2564 29648 2572
rect 29656 2564 29684 2572
rect 29692 2564 29712 2572
rect 29748 2572 29832 2592
rect 29748 2564 29768 2572
rect 29776 2564 29804 2572
rect 29812 2564 29832 2572
rect 29868 2572 29952 2592
rect 29868 2564 29888 2572
rect 29896 2564 29924 2572
rect 29932 2564 29952 2572
rect 29988 2572 30072 2592
rect 29988 2564 30008 2572
rect 30016 2564 30044 2572
rect 30052 2564 30072 2572
rect 30108 2572 30192 2592
rect 30108 2564 30128 2572
rect 30136 2564 30164 2572
rect 30172 2564 30192 2572
rect 30228 2572 30312 2592
rect 30228 2564 30248 2572
rect 30256 2564 30284 2572
rect 30292 2564 30312 2572
rect 30348 2572 30432 2592
rect 30348 2564 30368 2572
rect 30376 2564 30404 2572
rect 30412 2564 30432 2572
rect 30468 2572 30552 2592
rect 30468 2564 30488 2572
rect 30496 2564 30524 2572
rect 30532 2564 30552 2572
rect 30588 2572 30672 2592
rect 30588 2564 30608 2572
rect 30616 2564 30644 2572
rect 30652 2564 30672 2572
rect 30708 2572 30792 2592
rect 30708 2564 30728 2572
rect 30736 2564 30764 2572
rect 30772 2564 30792 2572
rect 30828 2572 30912 2592
rect 30828 2564 30848 2572
rect 30856 2564 30884 2572
rect 30892 2564 30912 2572
rect 30948 2572 31032 2592
rect 30948 2564 30968 2572
rect 30976 2564 31004 2572
rect 31012 2564 31032 2572
rect 31068 2572 31152 2592
rect 31068 2564 31088 2572
rect 31096 2564 31124 2572
rect 31132 2564 31152 2572
rect 31188 2572 31272 2592
rect 31188 2564 31208 2572
rect 31216 2564 31244 2572
rect 31252 2564 31272 2572
rect 31308 2572 31392 2592
rect 31308 2564 31328 2572
rect 31336 2564 31364 2572
rect 31372 2564 31392 2572
rect 31428 2572 31512 2592
rect 31428 2564 31448 2572
rect 31456 2564 31484 2572
rect 31492 2564 31512 2572
rect 31548 2572 31632 2592
rect 31548 2564 31568 2572
rect 31576 2564 31604 2572
rect 31612 2564 31632 2572
rect 31668 2572 31752 2592
rect 31668 2564 31688 2572
rect 31696 2564 31724 2572
rect 31732 2564 31752 2572
rect 31788 2572 31872 2592
rect 31788 2564 31808 2572
rect 31816 2564 31844 2572
rect 31852 2564 31872 2572
rect 31908 2572 31992 2592
rect 31908 2564 31928 2572
rect 31936 2564 31964 2572
rect 31972 2564 31992 2572
rect 32028 2572 32112 2592
rect 32028 2564 32048 2572
rect 32056 2564 32084 2572
rect 32092 2564 32112 2572
rect 32148 2572 32232 2592
rect 32148 2564 32168 2572
rect 32176 2564 32204 2572
rect 32212 2564 32232 2572
rect 32268 2572 32352 2592
rect 32268 2564 32288 2572
rect 32296 2564 32324 2572
rect 32332 2564 32352 2572
rect 32388 2572 32472 2592
rect 32388 2564 32408 2572
rect 32416 2564 32444 2572
rect 32452 2564 32472 2572
rect 32508 2572 32592 2592
rect 32508 2564 32528 2572
rect 32536 2564 32564 2572
rect 32572 2564 32592 2572
rect 32628 2572 32712 2592
rect 32628 2564 32648 2572
rect 32656 2564 32684 2572
rect 32692 2564 32712 2572
rect 32748 2572 32832 2592
rect 32748 2564 32768 2572
rect 32776 2564 32804 2572
rect 32812 2564 32832 2572
rect 32868 2572 32952 2592
rect 32868 2564 32888 2572
rect 32896 2564 32924 2572
rect 32932 2564 32952 2572
rect 32988 2572 33072 2592
rect 32988 2564 33008 2572
rect 33016 2564 33044 2572
rect 33052 2564 33072 2572
rect 33108 2572 33192 2592
rect 33108 2564 33128 2572
rect 33136 2564 33164 2572
rect 33172 2564 33192 2572
rect 33228 2572 33312 2592
rect 33228 2564 33248 2572
rect 33256 2564 33284 2572
rect 33292 2564 33312 2572
rect 33348 2572 33432 2592
rect 33348 2564 33368 2572
rect 33376 2564 33404 2572
rect 33412 2564 33432 2572
rect 33468 2572 33552 2592
rect 33468 2564 33488 2572
rect 33496 2564 33524 2572
rect 33532 2564 33552 2572
rect 33588 2572 33672 2592
rect 33588 2564 33608 2572
rect 33616 2564 33644 2572
rect 33652 2564 33672 2572
rect 33708 2572 33792 2592
rect 33708 2564 33728 2572
rect 33736 2564 33764 2572
rect 33772 2564 33792 2572
rect 33828 2572 33912 2592
rect 33828 2564 33848 2572
rect 33856 2564 33884 2572
rect 33892 2564 33912 2572
rect 33948 2572 34032 2592
rect 33948 2564 33968 2572
rect 33976 2564 34004 2572
rect 34012 2564 34032 2572
rect 34068 2572 34152 2592
rect 34068 2564 34088 2572
rect 34096 2564 34124 2572
rect 34132 2564 34152 2572
rect 34188 2572 34272 2592
rect 34188 2564 34208 2572
rect 34216 2564 34244 2572
rect 34252 2564 34272 2572
rect 34308 2572 34392 2592
rect 34308 2564 34328 2572
rect 34336 2564 34364 2572
rect 34372 2564 34392 2572
rect 34428 2572 34512 2592
rect 34428 2564 34448 2572
rect 34456 2564 34484 2572
rect 34492 2564 34512 2572
rect 34548 2572 34632 2592
rect 34548 2564 34568 2572
rect 34576 2564 34604 2572
rect 34612 2564 34632 2572
rect 34668 2572 34752 2592
rect 34668 2564 34688 2572
rect 34696 2564 34724 2572
rect 34732 2564 34752 2572
rect 34788 2572 34872 2592
rect 34788 2564 34808 2572
rect 34816 2564 34844 2572
rect 34852 2564 34872 2572
rect 34908 2572 34992 2592
rect 34908 2564 34928 2572
rect 34936 2564 34964 2572
rect 34972 2564 34992 2572
rect 35028 2572 35112 2592
rect 35028 2564 35048 2572
rect 35056 2564 35084 2572
rect 35092 2564 35112 2572
rect 35148 2572 35232 2592
rect 35148 2564 35168 2572
rect 35176 2564 35204 2572
rect 35212 2564 35232 2572
rect 35268 2572 35352 2592
rect 35268 2564 35288 2572
rect 35296 2564 35324 2572
rect 35332 2564 35352 2572
rect 35388 2572 35472 2592
rect 35388 2564 35408 2572
rect 35416 2564 35444 2572
rect 35452 2564 35472 2572
rect 35508 2572 35592 2592
rect 35508 2564 35528 2572
rect 35536 2564 35564 2572
rect 35572 2564 35592 2572
rect 35628 2572 35712 2592
rect 35628 2564 35648 2572
rect 35656 2564 35684 2572
rect 35692 2564 35712 2572
rect 35748 2572 35832 2592
rect 35748 2564 35768 2572
rect 35776 2564 35804 2572
rect 35812 2564 35832 2572
rect 35868 2572 35952 2592
rect 35868 2564 35888 2572
rect 35896 2564 35924 2572
rect 35932 2564 35952 2572
rect 35988 2572 36072 2592
rect 35988 2564 36008 2572
rect 36016 2564 36044 2572
rect 36052 2564 36072 2572
rect 36108 2572 36192 2592
rect 36108 2564 36128 2572
rect 36136 2564 36164 2572
rect 36172 2564 36192 2572
rect 36228 2572 36312 2592
rect 36228 2564 36248 2572
rect 36256 2564 36284 2572
rect 36292 2564 36312 2572
rect 36348 2572 36432 2592
rect 36348 2564 36368 2572
rect 36376 2564 36404 2572
rect 36412 2564 36432 2572
rect 36468 2572 36552 2592
rect 36468 2564 36488 2572
rect 36496 2564 36524 2572
rect 36532 2564 36552 2572
rect 36588 2572 36672 2592
rect 36588 2564 36608 2572
rect 36616 2564 36644 2572
rect 36652 2564 36672 2572
rect 36708 2572 36792 2592
rect 36708 2564 36728 2572
rect 36736 2564 36764 2572
rect 36772 2564 36792 2572
rect 36828 2572 36912 2592
rect 36828 2564 36848 2572
rect 36856 2564 36884 2572
rect 36892 2564 36912 2572
rect 36948 2572 37032 2592
rect 36948 2564 36968 2572
rect 36976 2564 37004 2572
rect 37012 2564 37032 2572
rect 37068 2572 37152 2592
rect 37068 2564 37088 2572
rect 37096 2564 37124 2572
rect 37132 2564 37152 2572
rect 37188 2572 37272 2592
rect 37188 2564 37208 2572
rect 37216 2564 37244 2572
rect 37252 2564 37272 2572
rect 37308 2572 37392 2592
rect 37308 2564 37328 2572
rect 37336 2564 37364 2572
rect 37372 2564 37392 2572
rect 37428 2572 37512 2592
rect 37428 2564 37448 2572
rect 37456 2564 37484 2572
rect 37492 2564 37512 2572
rect 37548 2572 37632 2592
rect 37548 2564 37568 2572
rect 37576 2564 37604 2572
rect 37612 2564 37632 2572
rect 37668 2572 37752 2592
rect 37668 2564 37688 2572
rect 37696 2564 37724 2572
rect 37732 2564 37752 2572
rect 37788 2572 37872 2592
rect 37788 2564 37808 2572
rect 37816 2564 37844 2572
rect 37852 2564 37872 2572
rect 37908 2572 37992 2592
rect 37908 2564 37928 2572
rect 37936 2564 37964 2572
rect 37972 2564 37992 2572
rect 38028 2572 38112 2592
rect 38028 2564 38048 2572
rect 38056 2564 38084 2572
rect 38092 2564 38112 2572
rect 38148 2572 38232 2592
rect 38148 2564 38168 2572
rect 38176 2564 38204 2572
rect 38212 2564 38232 2572
rect 38268 2572 38352 2592
rect 38268 2564 38288 2572
rect 38296 2564 38324 2572
rect 38332 2564 38352 2572
rect 38388 2572 38472 2592
rect 38388 2564 38408 2572
rect 38416 2564 38444 2572
rect 38452 2564 38472 2572
rect 38508 2572 38592 2592
rect 38508 2564 38528 2572
rect 38536 2564 38564 2572
rect 38572 2564 38592 2572
rect 38628 2572 38712 2592
rect 38628 2564 38648 2572
rect 38656 2564 38684 2572
rect 38692 2564 38712 2572
rect 38748 2572 38832 2592
rect 38748 2564 38768 2572
rect 38776 2564 38804 2572
rect 38812 2564 38832 2572
rect 38868 2572 38952 2592
rect 38868 2564 38888 2572
rect 38896 2564 38924 2572
rect 38932 2564 38952 2572
rect 38988 2572 39072 2592
rect 38988 2564 39008 2572
rect 39016 2564 39044 2572
rect 39052 2564 39072 2572
rect 39108 2572 39192 2592
rect 39108 2564 39128 2572
rect 39136 2564 39164 2572
rect 39172 2564 39192 2572
rect 39228 2572 39312 2592
rect 39228 2564 39248 2572
rect 39256 2564 39284 2572
rect 39292 2564 39312 2572
rect 39348 2572 39432 2592
rect 39348 2564 39368 2572
rect 39376 2564 39404 2572
rect 39412 2564 39432 2572
rect 39468 2572 39552 2592
rect 39468 2564 39488 2572
rect 39496 2564 39524 2572
rect 39532 2564 39552 2572
rect 39588 2572 39672 2592
rect 39588 2564 39608 2572
rect 39616 2564 39644 2572
rect 39652 2564 39672 2572
rect 39708 2572 39792 2592
rect 39708 2564 39728 2572
rect 39736 2564 39764 2572
rect 39772 2564 39792 2572
rect 39828 2572 39912 2592
rect 39828 2564 39848 2572
rect 39856 2564 39884 2572
rect 39892 2564 39912 2572
rect 39948 2572 40032 2592
rect 39948 2564 39968 2572
rect 39976 2564 40004 2572
rect 40012 2564 40032 2572
rect 40068 2572 40152 2592
rect 40068 2564 40088 2572
rect 40096 2564 40124 2572
rect 40132 2564 40152 2572
rect 40188 2572 40272 2592
rect 40188 2564 40208 2572
rect 40216 2564 40244 2572
rect 40252 2564 40272 2572
rect 40308 2572 40392 2592
rect 40308 2564 40328 2572
rect 40336 2564 40364 2572
rect 40372 2564 40392 2572
rect 40428 2572 40512 2592
rect 40428 2564 40448 2572
rect 40456 2564 40484 2572
rect 40492 2564 40512 2572
rect 40548 2572 40632 2592
rect 40548 2564 40568 2572
rect 40576 2564 40604 2572
rect 40612 2564 40632 2572
rect 40668 2572 40752 2592
rect 40668 2564 40688 2572
rect 40696 2564 40724 2572
rect 40732 2564 40752 2572
rect 40788 2572 40872 2592
rect 40788 2564 40808 2572
rect 40816 2564 40844 2572
rect 40852 2564 40872 2572
rect 40908 2572 40992 2592
rect 40908 2564 40928 2572
rect 40936 2564 40964 2572
rect 40972 2564 40992 2572
rect 41028 2572 41112 2592
rect 41028 2564 41048 2572
rect 41056 2564 41084 2572
rect 41092 2564 41112 2572
rect 41148 2572 41232 2592
rect 41148 2564 41168 2572
rect 41176 2564 41204 2572
rect 41212 2564 41232 2572
rect 41268 2572 41352 2592
rect 41268 2564 41288 2572
rect 41296 2564 41324 2572
rect 41332 2564 41352 2572
rect 41388 2572 41472 2592
rect 41388 2564 41408 2572
rect 41416 2564 41444 2572
rect 41452 2564 41472 2572
rect 41508 2572 41592 2592
rect 41508 2564 41528 2572
rect 41536 2564 41564 2572
rect 41572 2564 41592 2572
rect 41628 2572 41712 2592
rect 41628 2564 41648 2572
rect 41656 2564 41684 2572
rect 41692 2564 41712 2572
rect 41748 2572 41832 2592
rect 41748 2564 41768 2572
rect 41776 2564 41804 2572
rect 41812 2564 41832 2572
rect 41868 2572 41952 2592
rect 41868 2564 41888 2572
rect 41896 2564 41924 2572
rect 41932 2564 41952 2572
rect 41988 2572 42072 2592
rect 41988 2564 42008 2572
rect 42016 2564 42044 2572
rect 42052 2564 42072 2572
rect 42108 2572 42192 2592
rect 42108 2564 42128 2572
rect 42136 2564 42164 2572
rect 42172 2564 42192 2572
rect 42228 2572 42312 2592
rect 42228 2564 42248 2572
rect 42256 2564 42284 2572
rect 42292 2564 42312 2572
rect 42348 2572 42432 2592
rect 42348 2564 42368 2572
rect 42376 2564 42404 2572
rect 42412 2564 42432 2572
rect 42468 2572 42552 2592
rect 42468 2564 42488 2572
rect 42496 2564 42524 2572
rect 42532 2564 42552 2572
rect 42588 2572 42672 2592
rect 42588 2564 42608 2572
rect 42616 2564 42644 2572
rect 42652 2564 42672 2572
rect 42708 2572 42792 2592
rect 42708 2564 42728 2572
rect 42736 2564 42764 2572
rect 42772 2564 42792 2572
rect 42828 2572 42912 2592
rect 42828 2564 42848 2572
rect 42856 2564 42884 2572
rect 42892 2564 42912 2572
rect 42948 2572 43032 2592
rect 42948 2564 42968 2572
rect 42976 2564 43004 2572
rect 43012 2564 43032 2572
rect 43068 2572 43152 2592
rect 43068 2564 43088 2572
rect 43096 2564 43124 2572
rect 43132 2564 43152 2572
rect 43188 2572 43272 2592
rect 43188 2564 43208 2572
rect 43216 2564 43244 2572
rect 43252 2564 43272 2572
rect 43308 2572 43392 2592
rect 43308 2564 43328 2572
rect 43336 2564 43364 2572
rect 43372 2564 43392 2572
rect 43428 2572 43512 2592
rect 43428 2564 43448 2572
rect 43456 2564 43484 2572
rect 43492 2564 43512 2572
rect 43548 2572 43632 2592
rect 43548 2564 43568 2572
rect 43576 2564 43604 2572
rect 43612 2564 43632 2572
rect 43668 2572 43752 2592
rect 43668 2564 43688 2572
rect 43696 2564 43724 2572
rect 43732 2564 43752 2572
rect 43788 2572 43872 2592
rect 43788 2564 43808 2572
rect 43816 2564 43844 2572
rect 43852 2564 43872 2572
rect 43908 2572 43992 2592
rect 43908 2564 43928 2572
rect 43936 2564 43964 2572
rect 43972 2564 43992 2572
rect 44028 2572 44112 2592
rect 44028 2564 44048 2572
rect 44056 2564 44084 2572
rect 44092 2564 44112 2572
rect 44148 2572 44232 2592
rect 44148 2564 44168 2572
rect 44176 2564 44204 2572
rect 44212 2564 44232 2572
rect 44268 2572 44352 2592
rect 44268 2564 44288 2572
rect 44296 2564 44324 2572
rect 44332 2564 44352 2572
rect 44388 2572 44472 2592
rect 44388 2564 44408 2572
rect 44416 2564 44444 2572
rect 44452 2564 44472 2572
rect 44508 2572 44592 2592
rect 44508 2564 44528 2572
rect 44536 2564 44564 2572
rect 44572 2564 44592 2572
rect 44628 2572 44712 2592
rect 44628 2564 44648 2572
rect 44656 2564 44684 2572
rect 44692 2564 44712 2572
rect 44748 2572 44832 2592
rect 44748 2564 44768 2572
rect 44776 2564 44804 2572
rect 44812 2564 44832 2572
rect 44868 2572 44952 2592
rect 44868 2564 44888 2572
rect 44896 2564 44924 2572
rect 44932 2564 44952 2572
rect 44988 2572 45072 2592
rect 44988 2564 45008 2572
rect 45016 2564 45044 2572
rect 45052 2564 45072 2572
rect 45108 2572 45192 2592
rect 45108 2564 45128 2572
rect 45136 2564 45164 2572
rect 45172 2564 45192 2572
rect 45228 2572 45312 2592
rect 45228 2564 45248 2572
rect 45256 2564 45284 2572
rect 45292 2564 45312 2572
rect 45348 2572 45432 2592
rect 45348 2564 45368 2572
rect 45376 2564 45404 2572
rect 45412 2564 45432 2572
rect 45468 2572 45552 2592
rect 45468 2564 45488 2572
rect 45496 2564 45524 2572
rect 45532 2564 45552 2572
rect 45588 2572 45672 2592
rect 45588 2564 45608 2572
rect 45616 2564 45644 2572
rect 45652 2564 45672 2572
rect 25936 2536 25992 2564
rect 26056 2536 26112 2564
rect 26176 2536 26232 2564
rect 26296 2536 26352 2564
rect 26416 2536 26472 2564
rect 26536 2536 26592 2564
rect 26656 2536 26712 2564
rect 26776 2536 26832 2564
rect 26896 2536 26952 2564
rect 27016 2536 27072 2564
rect 27136 2536 27192 2564
rect 27256 2536 27312 2564
rect 27376 2536 27432 2564
rect 27496 2536 27552 2564
rect 27616 2536 27672 2564
rect 27736 2536 27792 2564
rect 27856 2536 27912 2564
rect 27976 2536 28032 2564
rect 28096 2536 28152 2564
rect 28216 2536 28272 2564
rect 28336 2536 28392 2564
rect 28456 2536 28512 2564
rect 28576 2536 28632 2564
rect 28696 2536 28752 2564
rect 28816 2536 28872 2564
rect 28936 2536 28992 2564
rect 29056 2536 29112 2564
rect 29176 2536 29232 2564
rect 29296 2536 29352 2564
rect 29416 2536 29472 2564
rect 29536 2536 29592 2564
rect 29656 2536 29712 2564
rect 29776 2536 29832 2564
rect 29896 2536 29952 2564
rect 30016 2536 30072 2564
rect 30136 2536 30192 2564
rect 30256 2536 30312 2564
rect 30376 2536 30432 2564
rect 30496 2536 30552 2564
rect 30616 2536 30672 2564
rect 30736 2536 30792 2564
rect 30856 2536 30912 2564
rect 30976 2536 31032 2564
rect 31096 2536 31152 2564
rect 31216 2536 31272 2564
rect 31336 2536 31392 2564
rect 31456 2536 31512 2564
rect 31576 2536 31632 2564
rect 31696 2536 31752 2564
rect 31816 2536 31872 2564
rect 31936 2536 31992 2564
rect 32056 2536 32112 2564
rect 32176 2536 32232 2564
rect 32296 2536 32352 2564
rect 32416 2536 32472 2564
rect 32536 2536 32592 2564
rect 32656 2536 32712 2564
rect 32776 2536 32832 2564
rect 32896 2536 32952 2564
rect 33016 2536 33072 2564
rect 33136 2536 33192 2564
rect 33256 2536 33312 2564
rect 33376 2536 33432 2564
rect 33496 2536 33552 2564
rect 33616 2536 33672 2564
rect 33736 2536 33792 2564
rect 33856 2536 33912 2564
rect 33976 2536 34032 2564
rect 34096 2536 34152 2564
rect 34216 2536 34272 2564
rect 34336 2536 34392 2564
rect 34456 2536 34512 2564
rect 34576 2536 34632 2564
rect 34696 2536 34752 2564
rect 34816 2536 34872 2564
rect 34936 2536 34992 2564
rect 35056 2536 35112 2564
rect 35176 2536 35232 2564
rect 35296 2536 35352 2564
rect 35416 2536 35472 2564
rect 35536 2536 35592 2564
rect 35656 2536 35712 2564
rect 35776 2536 35832 2564
rect 35896 2536 35952 2564
rect 36016 2536 36072 2564
rect 36136 2536 36192 2564
rect 36256 2536 36312 2564
rect 36376 2536 36432 2564
rect 36496 2536 36552 2564
rect 36616 2536 36672 2564
rect 36736 2536 36792 2564
rect 36856 2536 36912 2564
rect 36976 2536 37032 2564
rect 37096 2536 37152 2564
rect 37216 2536 37272 2564
rect 37336 2536 37392 2564
rect 37456 2536 37512 2564
rect 37576 2536 37632 2564
rect 37696 2536 37752 2564
rect 37816 2536 37872 2564
rect 37936 2536 37992 2564
rect 38056 2536 38112 2564
rect 38176 2536 38232 2564
rect 38296 2536 38352 2564
rect 38416 2536 38472 2564
rect 38536 2536 38592 2564
rect 38656 2536 38712 2564
rect 38776 2536 38832 2564
rect 38896 2536 38952 2564
rect 39016 2536 39072 2564
rect 39136 2536 39192 2564
rect 39256 2536 39312 2564
rect 39376 2536 39432 2564
rect 39496 2536 39552 2564
rect 39616 2536 39672 2564
rect 39736 2536 39792 2564
rect 39856 2536 39912 2564
rect 39976 2536 40032 2564
rect 40096 2536 40152 2564
rect 40216 2536 40272 2564
rect 40336 2536 40392 2564
rect 40456 2536 40512 2564
rect 40576 2536 40632 2564
rect 40696 2536 40752 2564
rect 40816 2536 40872 2564
rect 40936 2536 40992 2564
rect 41056 2536 41112 2564
rect 41176 2536 41232 2564
rect 41296 2536 41352 2564
rect 41416 2536 41472 2564
rect 41536 2536 41592 2564
rect 41656 2536 41712 2564
rect 41776 2536 41832 2564
rect 41896 2536 41952 2564
rect 42016 2536 42072 2564
rect 42136 2536 42192 2564
rect 42256 2536 42312 2564
rect 42376 2536 42432 2564
rect 42496 2536 42552 2564
rect 42616 2536 42672 2564
rect 42736 2536 42792 2564
rect 42856 2536 42912 2564
rect 42976 2536 43032 2564
rect 43096 2536 43152 2564
rect 43216 2536 43272 2564
rect 43336 2536 43392 2564
rect 43456 2536 43512 2564
rect 43576 2536 43632 2564
rect 43696 2536 43752 2564
rect 43816 2536 43872 2564
rect 43936 2536 43992 2564
rect 44056 2536 44112 2564
rect 44176 2536 44232 2564
rect 44296 2536 44352 2564
rect 44416 2536 44472 2564
rect 44536 2536 44592 2564
rect 44656 2536 44712 2564
rect 44776 2536 44832 2564
rect 44896 2536 44952 2564
rect 45016 2536 45072 2564
rect 45136 2536 45192 2564
rect 45256 2536 45312 2564
rect 45376 2536 45432 2564
rect 45496 2536 45552 2564
rect 45616 2536 45672 2564
rect 25848 1072 25932 1092
rect 25848 1064 25868 1072
rect 25876 1064 25904 1072
rect 25912 1064 25932 1072
rect 25968 1072 26052 1092
rect 25968 1064 25988 1072
rect 25996 1064 26024 1072
rect 26032 1064 26052 1072
rect 26088 1072 26172 1092
rect 26088 1064 26108 1072
rect 26116 1064 26144 1072
rect 26152 1064 26172 1072
rect 26208 1072 26292 1092
rect 26208 1064 26228 1072
rect 26236 1064 26264 1072
rect 26272 1064 26292 1072
rect 26328 1072 26412 1092
rect 26328 1064 26348 1072
rect 26356 1064 26384 1072
rect 26392 1064 26412 1072
rect 26448 1072 26532 1092
rect 26448 1064 26468 1072
rect 26476 1064 26504 1072
rect 26512 1064 26532 1072
rect 26568 1072 26652 1092
rect 26568 1064 26588 1072
rect 26596 1064 26624 1072
rect 26632 1064 26652 1072
rect 26688 1072 26772 1092
rect 26688 1064 26708 1072
rect 26716 1064 26744 1072
rect 26752 1064 26772 1072
rect 26808 1072 26892 1092
rect 26808 1064 26828 1072
rect 26836 1064 26864 1072
rect 26872 1064 26892 1072
rect 26928 1072 27012 1092
rect 26928 1064 26948 1072
rect 26956 1064 26984 1072
rect 26992 1064 27012 1072
rect 27048 1072 27132 1092
rect 27048 1064 27068 1072
rect 27076 1064 27104 1072
rect 27112 1064 27132 1072
rect 27168 1072 27252 1092
rect 27168 1064 27188 1072
rect 27196 1064 27224 1072
rect 27232 1064 27252 1072
rect 27288 1072 27372 1092
rect 27288 1064 27308 1072
rect 27316 1064 27344 1072
rect 27352 1064 27372 1072
rect 27408 1072 27492 1092
rect 27408 1064 27428 1072
rect 27436 1064 27464 1072
rect 27472 1064 27492 1072
rect 27528 1072 27612 1092
rect 27528 1064 27548 1072
rect 27556 1064 27584 1072
rect 27592 1064 27612 1072
rect 27648 1072 27732 1092
rect 27648 1064 27668 1072
rect 27676 1064 27704 1072
rect 27712 1064 27732 1072
rect 27768 1072 27852 1092
rect 27768 1064 27788 1072
rect 27796 1064 27824 1072
rect 27832 1064 27852 1072
rect 27888 1072 27972 1092
rect 27888 1064 27908 1072
rect 27916 1064 27944 1072
rect 27952 1064 27972 1072
rect 28008 1072 28092 1092
rect 28008 1064 28028 1072
rect 28036 1064 28064 1072
rect 28072 1064 28092 1072
rect 28128 1072 28212 1092
rect 28128 1064 28148 1072
rect 28156 1064 28184 1072
rect 28192 1064 28212 1072
rect 28248 1072 28332 1092
rect 28248 1064 28268 1072
rect 28276 1064 28304 1072
rect 28312 1064 28332 1072
rect 28368 1072 28452 1092
rect 28368 1064 28388 1072
rect 28396 1064 28424 1072
rect 28432 1064 28452 1072
rect 28488 1072 28572 1092
rect 28488 1064 28508 1072
rect 28516 1064 28544 1072
rect 28552 1064 28572 1072
rect 28608 1072 28692 1092
rect 28608 1064 28628 1072
rect 28636 1064 28664 1072
rect 28672 1064 28692 1072
rect 28728 1072 28812 1092
rect 28728 1064 28748 1072
rect 28756 1064 28784 1072
rect 28792 1064 28812 1072
rect 28848 1072 28932 1092
rect 28848 1064 28868 1072
rect 28876 1064 28904 1072
rect 28912 1064 28932 1072
rect 28968 1072 29052 1092
rect 28968 1064 28988 1072
rect 28996 1064 29024 1072
rect 29032 1064 29052 1072
rect 29088 1072 29172 1092
rect 29088 1064 29108 1072
rect 29116 1064 29144 1072
rect 29152 1064 29172 1072
rect 29208 1072 29292 1092
rect 29208 1064 29228 1072
rect 29236 1064 29264 1072
rect 29272 1064 29292 1072
rect 29328 1072 29412 1092
rect 29328 1064 29348 1072
rect 29356 1064 29384 1072
rect 29392 1064 29412 1072
rect 29448 1072 29532 1092
rect 29448 1064 29468 1072
rect 29476 1064 29504 1072
rect 29512 1064 29532 1072
rect 29568 1072 29652 1092
rect 29568 1064 29588 1072
rect 29596 1064 29624 1072
rect 29632 1064 29652 1072
rect 29688 1072 29772 1092
rect 29688 1064 29708 1072
rect 29716 1064 29744 1072
rect 29752 1064 29772 1072
rect 29808 1072 29892 1092
rect 29808 1064 29828 1072
rect 29836 1064 29864 1072
rect 29872 1064 29892 1072
rect 29928 1072 30012 1092
rect 29928 1064 29948 1072
rect 29956 1064 29984 1072
rect 29992 1064 30012 1072
rect 30048 1072 30132 1092
rect 30048 1064 30068 1072
rect 30076 1064 30104 1072
rect 30112 1064 30132 1072
rect 30168 1072 30252 1092
rect 30168 1064 30188 1072
rect 30196 1064 30224 1072
rect 30232 1064 30252 1072
rect 30288 1072 30372 1092
rect 30288 1064 30308 1072
rect 30316 1064 30344 1072
rect 30352 1064 30372 1072
rect 30408 1072 30492 1092
rect 30408 1064 30428 1072
rect 30436 1064 30464 1072
rect 30472 1064 30492 1072
rect 30528 1072 30612 1092
rect 30528 1064 30548 1072
rect 30556 1064 30584 1072
rect 30592 1064 30612 1072
rect 30648 1072 30732 1092
rect 30648 1064 30668 1072
rect 30676 1064 30704 1072
rect 30712 1064 30732 1072
rect 30768 1072 30852 1092
rect 30768 1064 30788 1072
rect 30796 1064 30824 1072
rect 30832 1064 30852 1072
rect 30888 1072 30972 1092
rect 30888 1064 30908 1072
rect 30916 1064 30944 1072
rect 30952 1064 30972 1072
rect 31008 1072 31092 1092
rect 31008 1064 31028 1072
rect 31036 1064 31064 1072
rect 31072 1064 31092 1072
rect 31128 1072 31212 1092
rect 31128 1064 31148 1072
rect 31156 1064 31184 1072
rect 31192 1064 31212 1072
rect 31248 1072 31332 1092
rect 31248 1064 31268 1072
rect 31276 1064 31304 1072
rect 31312 1064 31332 1072
rect 31368 1072 31452 1092
rect 31368 1064 31388 1072
rect 31396 1064 31424 1072
rect 31432 1064 31452 1072
rect 31488 1072 31572 1092
rect 31488 1064 31508 1072
rect 31516 1064 31544 1072
rect 31552 1064 31572 1072
rect 31608 1072 31692 1092
rect 31608 1064 31628 1072
rect 31636 1064 31664 1072
rect 31672 1064 31692 1072
rect 31728 1072 31812 1092
rect 31728 1064 31748 1072
rect 31756 1064 31784 1072
rect 31792 1064 31812 1072
rect 31848 1072 31932 1092
rect 31848 1064 31868 1072
rect 31876 1064 31904 1072
rect 31912 1064 31932 1072
rect 31968 1072 32052 1092
rect 31968 1064 31988 1072
rect 31996 1064 32024 1072
rect 32032 1064 32052 1072
rect 32088 1072 32172 1092
rect 32088 1064 32108 1072
rect 32116 1064 32144 1072
rect 32152 1064 32172 1072
rect 32208 1072 32292 1092
rect 32208 1064 32228 1072
rect 32236 1064 32264 1072
rect 32272 1064 32292 1072
rect 32328 1072 32412 1092
rect 32328 1064 32348 1072
rect 32356 1064 32384 1072
rect 32392 1064 32412 1072
rect 32448 1072 32532 1092
rect 32448 1064 32468 1072
rect 32476 1064 32504 1072
rect 32512 1064 32532 1072
rect 32568 1072 32652 1092
rect 32568 1064 32588 1072
rect 32596 1064 32624 1072
rect 32632 1064 32652 1072
rect 32688 1072 32772 1092
rect 32688 1064 32708 1072
rect 32716 1064 32744 1072
rect 32752 1064 32772 1072
rect 32808 1072 32892 1092
rect 32808 1064 32828 1072
rect 32836 1064 32864 1072
rect 32872 1064 32892 1072
rect 32928 1072 33012 1092
rect 32928 1064 32948 1072
rect 32956 1064 32984 1072
rect 32992 1064 33012 1072
rect 33048 1072 33132 1092
rect 33048 1064 33068 1072
rect 33076 1064 33104 1072
rect 33112 1064 33132 1072
rect 33168 1072 33252 1092
rect 33168 1064 33188 1072
rect 33196 1064 33224 1072
rect 33232 1064 33252 1072
rect 33288 1072 33372 1092
rect 33288 1064 33308 1072
rect 33316 1064 33344 1072
rect 33352 1064 33372 1072
rect 33408 1072 33492 1092
rect 33408 1064 33428 1072
rect 33436 1064 33464 1072
rect 33472 1064 33492 1072
rect 33528 1072 33612 1092
rect 33528 1064 33548 1072
rect 33556 1064 33584 1072
rect 33592 1064 33612 1072
rect 33648 1072 33732 1092
rect 33648 1064 33668 1072
rect 33676 1064 33704 1072
rect 33712 1064 33732 1072
rect 33768 1072 33852 1092
rect 33768 1064 33788 1072
rect 33796 1064 33824 1072
rect 33832 1064 33852 1072
rect 33888 1072 33972 1092
rect 33888 1064 33908 1072
rect 33916 1064 33944 1072
rect 33952 1064 33972 1072
rect 34008 1072 34092 1092
rect 34008 1064 34028 1072
rect 34036 1064 34064 1072
rect 34072 1064 34092 1072
rect 34128 1072 34212 1092
rect 34128 1064 34148 1072
rect 34156 1064 34184 1072
rect 34192 1064 34212 1072
rect 34248 1072 34332 1092
rect 34248 1064 34268 1072
rect 34276 1064 34304 1072
rect 34312 1064 34332 1072
rect 34368 1072 34452 1092
rect 34368 1064 34388 1072
rect 34396 1064 34424 1072
rect 34432 1064 34452 1072
rect 34488 1072 34572 1092
rect 34488 1064 34508 1072
rect 34516 1064 34544 1072
rect 34552 1064 34572 1072
rect 34608 1072 34692 1092
rect 34608 1064 34628 1072
rect 34636 1064 34664 1072
rect 34672 1064 34692 1072
rect 34728 1072 34812 1092
rect 34728 1064 34748 1072
rect 34756 1064 34784 1072
rect 34792 1064 34812 1072
rect 34848 1072 34932 1092
rect 34848 1064 34868 1072
rect 34876 1064 34904 1072
rect 34912 1064 34932 1072
rect 34968 1072 35052 1092
rect 34968 1064 34988 1072
rect 34996 1064 35024 1072
rect 35032 1064 35052 1072
rect 35088 1072 35172 1092
rect 35088 1064 35108 1072
rect 35116 1064 35144 1072
rect 35152 1064 35172 1072
rect 35208 1072 35292 1092
rect 35208 1064 35228 1072
rect 35236 1064 35264 1072
rect 35272 1064 35292 1072
rect 35328 1072 35412 1092
rect 35328 1064 35348 1072
rect 35356 1064 35384 1072
rect 35392 1064 35412 1072
rect 35448 1072 35532 1092
rect 35448 1064 35468 1072
rect 35476 1064 35504 1072
rect 35512 1064 35532 1072
rect 35568 1072 35652 1092
rect 35568 1064 35588 1072
rect 35596 1064 35624 1072
rect 35632 1064 35652 1072
rect 35688 1072 35772 1092
rect 35688 1064 35708 1072
rect 35716 1064 35744 1072
rect 35752 1064 35772 1072
rect 35808 1072 35892 1092
rect 35808 1064 35828 1072
rect 35836 1064 35864 1072
rect 35872 1064 35892 1072
rect 35928 1072 36012 1092
rect 35928 1064 35948 1072
rect 35956 1064 35984 1072
rect 35992 1064 36012 1072
rect 36048 1072 36132 1092
rect 36048 1064 36068 1072
rect 36076 1064 36104 1072
rect 36112 1064 36132 1072
rect 36168 1072 36252 1092
rect 36168 1064 36188 1072
rect 36196 1064 36224 1072
rect 36232 1064 36252 1072
rect 36288 1072 36372 1092
rect 36288 1064 36308 1072
rect 36316 1064 36344 1072
rect 36352 1064 36372 1072
rect 36408 1072 36492 1092
rect 36408 1064 36428 1072
rect 36436 1064 36464 1072
rect 36472 1064 36492 1072
rect 36528 1072 36612 1092
rect 36528 1064 36548 1072
rect 36556 1064 36584 1072
rect 36592 1064 36612 1072
rect 36648 1072 36732 1092
rect 36648 1064 36668 1072
rect 36676 1064 36704 1072
rect 36712 1064 36732 1072
rect 36768 1072 36852 1092
rect 36768 1064 36788 1072
rect 36796 1064 36824 1072
rect 36832 1064 36852 1072
rect 36888 1072 36972 1092
rect 36888 1064 36908 1072
rect 36916 1064 36944 1072
rect 36952 1064 36972 1072
rect 37008 1072 37092 1092
rect 37008 1064 37028 1072
rect 37036 1064 37064 1072
rect 37072 1064 37092 1072
rect 37128 1072 37212 1092
rect 37128 1064 37148 1072
rect 37156 1064 37184 1072
rect 37192 1064 37212 1072
rect 37248 1072 37332 1092
rect 37248 1064 37268 1072
rect 37276 1064 37304 1072
rect 37312 1064 37332 1072
rect 37368 1072 37452 1092
rect 37368 1064 37388 1072
rect 37396 1064 37424 1072
rect 37432 1064 37452 1072
rect 37488 1072 37572 1092
rect 37488 1064 37508 1072
rect 37516 1064 37544 1072
rect 37552 1064 37572 1072
rect 37608 1072 37692 1092
rect 37608 1064 37628 1072
rect 37636 1064 37664 1072
rect 37672 1064 37692 1072
rect 37728 1072 37812 1092
rect 37728 1064 37748 1072
rect 37756 1064 37784 1072
rect 37792 1064 37812 1072
rect 37848 1072 37932 1092
rect 37848 1064 37868 1072
rect 37876 1064 37904 1072
rect 37912 1064 37932 1072
rect 37968 1072 38052 1092
rect 37968 1064 37988 1072
rect 37996 1064 38024 1072
rect 38032 1064 38052 1072
rect 38088 1072 38172 1092
rect 38088 1064 38108 1072
rect 38116 1064 38144 1072
rect 38152 1064 38172 1072
rect 38208 1072 38292 1092
rect 38208 1064 38228 1072
rect 38236 1064 38264 1072
rect 38272 1064 38292 1072
rect 38328 1072 38412 1092
rect 38328 1064 38348 1072
rect 38356 1064 38384 1072
rect 38392 1064 38412 1072
rect 38448 1072 38532 1092
rect 38448 1064 38468 1072
rect 38476 1064 38504 1072
rect 38512 1064 38532 1072
rect 38568 1072 38652 1092
rect 38568 1064 38588 1072
rect 38596 1064 38624 1072
rect 38632 1064 38652 1072
rect 38688 1072 38772 1092
rect 38688 1064 38708 1072
rect 38716 1064 38744 1072
rect 38752 1064 38772 1072
rect 38808 1072 38892 1092
rect 38808 1064 38828 1072
rect 38836 1064 38864 1072
rect 38872 1064 38892 1072
rect 38928 1072 39012 1092
rect 38928 1064 38948 1072
rect 38956 1064 38984 1072
rect 38992 1064 39012 1072
rect 39048 1072 39132 1092
rect 39048 1064 39068 1072
rect 39076 1064 39104 1072
rect 39112 1064 39132 1072
rect 39168 1072 39252 1092
rect 39168 1064 39188 1072
rect 39196 1064 39224 1072
rect 39232 1064 39252 1072
rect 39288 1072 39372 1092
rect 39288 1064 39308 1072
rect 39316 1064 39344 1072
rect 39352 1064 39372 1072
rect 39408 1072 39492 1092
rect 39408 1064 39428 1072
rect 39436 1064 39464 1072
rect 39472 1064 39492 1072
rect 39528 1072 39612 1092
rect 39528 1064 39548 1072
rect 39556 1064 39584 1072
rect 39592 1064 39612 1072
rect 39648 1072 39732 1092
rect 39648 1064 39668 1072
rect 39676 1064 39704 1072
rect 39712 1064 39732 1072
rect 39768 1072 39852 1092
rect 39768 1064 39788 1072
rect 39796 1064 39824 1072
rect 39832 1064 39852 1072
rect 39888 1072 39972 1092
rect 39888 1064 39908 1072
rect 39916 1064 39944 1072
rect 39952 1064 39972 1072
rect 40008 1072 40092 1092
rect 40008 1064 40028 1072
rect 40036 1064 40064 1072
rect 40072 1064 40092 1072
rect 40128 1072 40212 1092
rect 40128 1064 40148 1072
rect 40156 1064 40184 1072
rect 40192 1064 40212 1072
rect 40248 1072 40332 1092
rect 40248 1064 40268 1072
rect 40276 1064 40304 1072
rect 40312 1064 40332 1072
rect 40368 1072 40452 1092
rect 40368 1064 40388 1072
rect 40396 1064 40424 1072
rect 40432 1064 40452 1072
rect 40488 1072 40572 1092
rect 40488 1064 40508 1072
rect 40516 1064 40544 1072
rect 40552 1064 40572 1072
rect 40608 1072 40692 1092
rect 40608 1064 40628 1072
rect 40636 1064 40664 1072
rect 40672 1064 40692 1072
rect 40728 1072 40812 1092
rect 40728 1064 40748 1072
rect 40756 1064 40784 1072
rect 40792 1064 40812 1072
rect 40848 1072 40932 1092
rect 40848 1064 40868 1072
rect 40876 1064 40904 1072
rect 40912 1064 40932 1072
rect 40968 1072 41052 1092
rect 40968 1064 40988 1072
rect 40996 1064 41024 1072
rect 41032 1064 41052 1072
rect 41088 1072 41172 1092
rect 41088 1064 41108 1072
rect 41116 1064 41144 1072
rect 41152 1064 41172 1072
rect 41208 1072 41292 1092
rect 41208 1064 41228 1072
rect 41236 1064 41264 1072
rect 41272 1064 41292 1072
rect 41328 1072 41412 1092
rect 41328 1064 41348 1072
rect 41356 1064 41384 1072
rect 41392 1064 41412 1072
rect 41448 1072 41532 1092
rect 41448 1064 41468 1072
rect 41476 1064 41504 1072
rect 41512 1064 41532 1072
rect 41568 1072 41652 1092
rect 41568 1064 41588 1072
rect 41596 1064 41624 1072
rect 41632 1064 41652 1072
rect 41688 1072 41772 1092
rect 41688 1064 41708 1072
rect 41716 1064 41744 1072
rect 41752 1064 41772 1072
rect 41808 1072 41892 1092
rect 41808 1064 41828 1072
rect 41836 1064 41864 1072
rect 41872 1064 41892 1072
rect 41928 1072 42012 1092
rect 41928 1064 41948 1072
rect 41956 1064 41984 1072
rect 41992 1064 42012 1072
rect 42048 1072 42132 1092
rect 42048 1064 42068 1072
rect 42076 1064 42104 1072
rect 42112 1064 42132 1072
rect 42168 1072 42252 1092
rect 42168 1064 42188 1072
rect 42196 1064 42224 1072
rect 42232 1064 42252 1072
rect 42288 1072 42372 1092
rect 42288 1064 42308 1072
rect 42316 1064 42344 1072
rect 42352 1064 42372 1072
rect 42408 1072 42492 1092
rect 42408 1064 42428 1072
rect 42436 1064 42464 1072
rect 42472 1064 42492 1072
rect 42528 1072 42612 1092
rect 42528 1064 42548 1072
rect 42556 1064 42584 1072
rect 42592 1064 42612 1072
rect 42648 1072 42732 1092
rect 42648 1064 42668 1072
rect 42676 1064 42704 1072
rect 42712 1064 42732 1072
rect 42768 1072 42852 1092
rect 42768 1064 42788 1072
rect 42796 1064 42824 1072
rect 42832 1064 42852 1072
rect 42888 1072 42972 1092
rect 42888 1064 42908 1072
rect 42916 1064 42944 1072
rect 42952 1064 42972 1072
rect 43008 1072 43092 1092
rect 43008 1064 43028 1072
rect 43036 1064 43064 1072
rect 43072 1064 43092 1072
rect 43128 1072 43212 1092
rect 43128 1064 43148 1072
rect 43156 1064 43184 1072
rect 43192 1064 43212 1072
rect 43248 1072 43332 1092
rect 43248 1064 43268 1072
rect 43276 1064 43304 1072
rect 43312 1064 43332 1072
rect 43368 1072 43452 1092
rect 43368 1064 43388 1072
rect 43396 1064 43424 1072
rect 43432 1064 43452 1072
rect 43488 1072 43572 1092
rect 43488 1064 43508 1072
rect 43516 1064 43544 1072
rect 43552 1064 43572 1072
rect 43608 1072 43692 1092
rect 43608 1064 43628 1072
rect 43636 1064 43664 1072
rect 43672 1064 43692 1072
rect 43728 1072 43812 1092
rect 43728 1064 43748 1072
rect 43756 1064 43784 1072
rect 43792 1064 43812 1072
rect 43848 1072 43932 1092
rect 43848 1064 43868 1072
rect 43876 1064 43904 1072
rect 43912 1064 43932 1072
rect 43968 1072 44052 1092
rect 43968 1064 43988 1072
rect 43996 1064 44024 1072
rect 44032 1064 44052 1072
rect 44088 1072 44172 1092
rect 44088 1064 44108 1072
rect 44116 1064 44144 1072
rect 44152 1064 44172 1072
rect 44208 1072 44292 1092
rect 44208 1064 44228 1072
rect 44236 1064 44264 1072
rect 44272 1064 44292 1072
rect 44328 1072 44412 1092
rect 44328 1064 44348 1072
rect 44356 1064 44384 1072
rect 44392 1064 44412 1072
rect 44448 1072 44532 1092
rect 44448 1064 44468 1072
rect 44476 1064 44504 1072
rect 44512 1064 44532 1072
rect 44568 1072 44652 1092
rect 44568 1064 44588 1072
rect 44596 1064 44624 1072
rect 44632 1064 44652 1072
rect 44688 1072 44772 1092
rect 44688 1064 44708 1072
rect 44716 1064 44744 1072
rect 44752 1064 44772 1072
rect 44808 1072 44892 1092
rect 44808 1064 44828 1072
rect 44836 1064 44864 1072
rect 44872 1064 44892 1072
rect 44928 1072 45012 1092
rect 44928 1064 44948 1072
rect 44956 1064 44984 1072
rect 44992 1064 45012 1072
rect 45048 1072 45132 1092
rect 45048 1064 45068 1072
rect 45076 1064 45104 1072
rect 45112 1064 45132 1072
rect 45168 1072 45252 1092
rect 45168 1064 45188 1072
rect 45196 1064 45224 1072
rect 45232 1064 45252 1072
rect 45288 1072 45372 1092
rect 45288 1064 45308 1072
rect 45316 1064 45344 1072
rect 45352 1064 45372 1072
rect 45408 1072 45492 1092
rect 45408 1064 45428 1072
rect 45436 1064 45464 1072
rect 45472 1064 45492 1072
rect 45528 1072 45612 1092
rect 45528 1064 45548 1072
rect 45556 1064 45584 1072
rect 45592 1064 45612 1072
rect 25876 1036 25932 1064
rect 25996 1036 26052 1064
rect 26116 1036 26172 1064
rect 26236 1036 26292 1064
rect 26356 1036 26412 1064
rect 26476 1036 26532 1064
rect 26596 1036 26652 1064
rect 26716 1036 26772 1064
rect 26836 1036 26892 1064
rect 26956 1036 27012 1064
rect 27076 1036 27132 1064
rect 27196 1036 27252 1064
rect 27316 1036 27372 1064
rect 27436 1036 27492 1064
rect 27556 1036 27612 1064
rect 27676 1036 27732 1064
rect 27796 1036 27852 1064
rect 27916 1036 27972 1064
rect 28036 1036 28092 1064
rect 28156 1036 28212 1064
rect 28276 1036 28332 1064
rect 28396 1036 28452 1064
rect 28516 1036 28572 1064
rect 28636 1036 28692 1064
rect 28756 1036 28812 1064
rect 28876 1036 28932 1064
rect 28996 1036 29052 1064
rect 29116 1036 29172 1064
rect 29236 1036 29292 1064
rect 29356 1036 29412 1064
rect 29476 1036 29532 1064
rect 29596 1036 29652 1064
rect 29716 1036 29772 1064
rect 29836 1036 29892 1064
rect 29956 1036 30012 1064
rect 30076 1036 30132 1064
rect 30196 1036 30252 1064
rect 30316 1036 30372 1064
rect 30436 1036 30492 1064
rect 30556 1036 30612 1064
rect 30676 1036 30732 1064
rect 30796 1036 30852 1064
rect 30916 1036 30972 1064
rect 31036 1036 31092 1064
rect 31156 1036 31212 1064
rect 31276 1036 31332 1064
rect 31396 1036 31452 1064
rect 31516 1036 31572 1064
rect 31636 1036 31692 1064
rect 31756 1036 31812 1064
rect 31876 1036 31932 1064
rect 31996 1036 32052 1064
rect 32116 1036 32172 1064
rect 32236 1036 32292 1064
rect 32356 1036 32412 1064
rect 32476 1036 32532 1064
rect 32596 1036 32652 1064
rect 32716 1036 32772 1064
rect 32836 1036 32892 1064
rect 32956 1036 33012 1064
rect 33076 1036 33132 1064
rect 33196 1036 33252 1064
rect 33316 1036 33372 1064
rect 33436 1036 33492 1064
rect 33556 1036 33612 1064
rect 33676 1036 33732 1064
rect 33796 1036 33852 1064
rect 33916 1036 33972 1064
rect 34036 1036 34092 1064
rect 34156 1036 34212 1064
rect 34276 1036 34332 1064
rect 34396 1036 34452 1064
rect 34516 1036 34572 1064
rect 34636 1036 34692 1064
rect 34756 1036 34812 1064
rect 34876 1036 34932 1064
rect 34996 1036 35052 1064
rect 35116 1036 35172 1064
rect 35236 1036 35292 1064
rect 35356 1036 35412 1064
rect 35476 1036 35532 1064
rect 35596 1036 35652 1064
rect 35716 1036 35772 1064
rect 35836 1036 35892 1064
rect 35956 1036 36012 1064
rect 36076 1036 36132 1064
rect 36196 1036 36252 1064
rect 36316 1036 36372 1064
rect 36436 1036 36492 1064
rect 36556 1036 36612 1064
rect 36676 1036 36732 1064
rect 36796 1036 36852 1064
rect 36916 1036 36972 1064
rect 37036 1036 37092 1064
rect 37156 1036 37212 1064
rect 37276 1036 37332 1064
rect 37396 1036 37452 1064
rect 37516 1036 37572 1064
rect 37636 1036 37692 1064
rect 37756 1036 37812 1064
rect 37876 1036 37932 1064
rect 37996 1036 38052 1064
rect 38116 1036 38172 1064
rect 38236 1036 38292 1064
rect 38356 1036 38412 1064
rect 38476 1036 38532 1064
rect 38596 1036 38652 1064
rect 38716 1036 38772 1064
rect 38836 1036 38892 1064
rect 38956 1036 39012 1064
rect 39076 1036 39132 1064
rect 39196 1036 39252 1064
rect 39316 1036 39372 1064
rect 39436 1036 39492 1064
rect 39556 1036 39612 1064
rect 39676 1036 39732 1064
rect 39796 1036 39852 1064
rect 39916 1036 39972 1064
rect 40036 1036 40092 1064
rect 40156 1036 40212 1064
rect 40276 1036 40332 1064
rect 40396 1036 40452 1064
rect 40516 1036 40572 1064
rect 40636 1036 40692 1064
rect 40756 1036 40812 1064
rect 40876 1036 40932 1064
rect 40996 1036 41052 1064
rect 41116 1036 41172 1064
rect 41236 1036 41292 1064
rect 41356 1036 41412 1064
rect 41476 1036 41532 1064
rect 41596 1036 41652 1064
rect 41716 1036 41772 1064
rect 41836 1036 41892 1064
rect 41956 1036 42012 1064
rect 42076 1036 42132 1064
rect 42196 1036 42252 1064
rect 42316 1036 42372 1064
rect 42436 1036 42492 1064
rect 42556 1036 42612 1064
rect 42676 1036 42732 1064
rect 42796 1036 42852 1064
rect 42916 1036 42972 1064
rect 43036 1036 43092 1064
rect 43156 1036 43212 1064
rect 43276 1036 43332 1064
rect 43396 1036 43452 1064
rect 43516 1036 43572 1064
rect 43636 1036 43692 1064
rect 43756 1036 43812 1064
rect 43876 1036 43932 1064
rect 43996 1036 44052 1064
rect 44116 1036 44172 1064
rect 44236 1036 44292 1064
rect 44356 1036 44412 1064
rect 44476 1036 44532 1064
rect 44596 1036 44652 1064
rect 44716 1036 44772 1064
rect 44836 1036 44892 1064
rect 44956 1036 45012 1064
rect 45076 1036 45132 1064
rect 45196 1036 45252 1064
rect 45316 1036 45372 1064
rect 45436 1036 45492 1064
rect 45556 1036 45612 1064
rect 25848 892 25932 912
rect 25848 884 25868 892
rect 25876 884 25904 892
rect 25912 884 25932 892
rect 25968 892 26052 912
rect 25968 884 25988 892
rect 25996 884 26024 892
rect 26032 884 26052 892
rect 26088 892 26172 912
rect 26088 884 26108 892
rect 26116 884 26144 892
rect 26152 884 26172 892
rect 26208 892 26292 912
rect 26208 884 26228 892
rect 26236 884 26264 892
rect 26272 884 26292 892
rect 26328 892 26412 912
rect 26328 884 26348 892
rect 26356 884 26384 892
rect 26392 884 26412 892
rect 26448 892 26532 912
rect 26448 884 26468 892
rect 26476 884 26504 892
rect 26512 884 26532 892
rect 26568 892 26652 912
rect 26568 884 26588 892
rect 26596 884 26624 892
rect 26632 884 26652 892
rect 26688 892 26772 912
rect 26688 884 26708 892
rect 26716 884 26744 892
rect 26752 884 26772 892
rect 26808 892 26892 912
rect 26808 884 26828 892
rect 26836 884 26864 892
rect 26872 884 26892 892
rect 26928 892 27012 912
rect 26928 884 26948 892
rect 26956 884 26984 892
rect 26992 884 27012 892
rect 27048 892 27132 912
rect 27048 884 27068 892
rect 27076 884 27104 892
rect 27112 884 27132 892
rect 27168 892 27252 912
rect 27168 884 27188 892
rect 27196 884 27224 892
rect 27232 884 27252 892
rect 27288 892 27372 912
rect 27288 884 27308 892
rect 27316 884 27344 892
rect 27352 884 27372 892
rect 27408 892 27492 912
rect 27408 884 27428 892
rect 27436 884 27464 892
rect 27472 884 27492 892
rect 27528 892 27612 912
rect 27528 884 27548 892
rect 27556 884 27584 892
rect 27592 884 27612 892
rect 27648 892 27732 912
rect 27648 884 27668 892
rect 27676 884 27704 892
rect 27712 884 27732 892
rect 27768 892 27852 912
rect 27768 884 27788 892
rect 27796 884 27824 892
rect 27832 884 27852 892
rect 27888 892 27972 912
rect 27888 884 27908 892
rect 27916 884 27944 892
rect 27952 884 27972 892
rect 28008 892 28092 912
rect 28008 884 28028 892
rect 28036 884 28064 892
rect 28072 884 28092 892
rect 28128 892 28212 912
rect 28128 884 28148 892
rect 28156 884 28184 892
rect 28192 884 28212 892
rect 28248 892 28332 912
rect 28248 884 28268 892
rect 28276 884 28304 892
rect 28312 884 28332 892
rect 28368 892 28452 912
rect 28368 884 28388 892
rect 28396 884 28424 892
rect 28432 884 28452 892
rect 28488 892 28572 912
rect 28488 884 28508 892
rect 28516 884 28544 892
rect 28552 884 28572 892
rect 28608 892 28692 912
rect 28608 884 28628 892
rect 28636 884 28664 892
rect 28672 884 28692 892
rect 28728 892 28812 912
rect 28728 884 28748 892
rect 28756 884 28784 892
rect 28792 884 28812 892
rect 28848 892 28932 912
rect 28848 884 28868 892
rect 28876 884 28904 892
rect 28912 884 28932 892
rect 28968 892 29052 912
rect 28968 884 28988 892
rect 28996 884 29024 892
rect 29032 884 29052 892
rect 29088 892 29172 912
rect 29088 884 29108 892
rect 29116 884 29144 892
rect 29152 884 29172 892
rect 29208 892 29292 912
rect 29208 884 29228 892
rect 29236 884 29264 892
rect 29272 884 29292 892
rect 29328 892 29412 912
rect 29328 884 29348 892
rect 29356 884 29384 892
rect 29392 884 29412 892
rect 29448 892 29532 912
rect 29448 884 29468 892
rect 29476 884 29504 892
rect 29512 884 29532 892
rect 29568 892 29652 912
rect 29568 884 29588 892
rect 29596 884 29624 892
rect 29632 884 29652 892
rect 29688 892 29772 912
rect 29688 884 29708 892
rect 29716 884 29744 892
rect 29752 884 29772 892
rect 29808 892 29892 912
rect 29808 884 29828 892
rect 29836 884 29864 892
rect 29872 884 29892 892
rect 29928 892 30012 912
rect 29928 884 29948 892
rect 29956 884 29984 892
rect 29992 884 30012 892
rect 30048 892 30132 912
rect 30048 884 30068 892
rect 30076 884 30104 892
rect 30112 884 30132 892
rect 30168 892 30252 912
rect 30168 884 30188 892
rect 30196 884 30224 892
rect 30232 884 30252 892
rect 30288 892 30372 912
rect 30288 884 30308 892
rect 30316 884 30344 892
rect 30352 884 30372 892
rect 30408 892 30492 912
rect 30408 884 30428 892
rect 30436 884 30464 892
rect 30472 884 30492 892
rect 30528 892 30612 912
rect 30528 884 30548 892
rect 30556 884 30584 892
rect 30592 884 30612 892
rect 30648 892 30732 912
rect 30648 884 30668 892
rect 30676 884 30704 892
rect 30712 884 30732 892
rect 30768 892 30852 912
rect 30768 884 30788 892
rect 30796 884 30824 892
rect 30832 884 30852 892
rect 30888 892 30972 912
rect 30888 884 30908 892
rect 30916 884 30944 892
rect 30952 884 30972 892
rect 31008 892 31092 912
rect 31008 884 31028 892
rect 31036 884 31064 892
rect 31072 884 31092 892
rect 31128 892 31212 912
rect 31128 884 31148 892
rect 31156 884 31184 892
rect 31192 884 31212 892
rect 31248 892 31332 912
rect 31248 884 31268 892
rect 31276 884 31304 892
rect 31312 884 31332 892
rect 31368 892 31452 912
rect 31368 884 31388 892
rect 31396 884 31424 892
rect 31432 884 31452 892
rect 31488 892 31572 912
rect 31488 884 31508 892
rect 31516 884 31544 892
rect 31552 884 31572 892
rect 31608 892 31692 912
rect 31608 884 31628 892
rect 31636 884 31664 892
rect 31672 884 31692 892
rect 31728 892 31812 912
rect 31728 884 31748 892
rect 31756 884 31784 892
rect 31792 884 31812 892
rect 31848 892 31932 912
rect 31848 884 31868 892
rect 31876 884 31904 892
rect 31912 884 31932 892
rect 31968 892 32052 912
rect 31968 884 31988 892
rect 31996 884 32024 892
rect 32032 884 32052 892
rect 32088 892 32172 912
rect 32088 884 32108 892
rect 32116 884 32144 892
rect 32152 884 32172 892
rect 32208 892 32292 912
rect 32208 884 32228 892
rect 32236 884 32264 892
rect 32272 884 32292 892
rect 32328 892 32412 912
rect 32328 884 32348 892
rect 32356 884 32384 892
rect 32392 884 32412 892
rect 32448 892 32532 912
rect 32448 884 32468 892
rect 32476 884 32504 892
rect 32512 884 32532 892
rect 32568 892 32652 912
rect 32568 884 32588 892
rect 32596 884 32624 892
rect 32632 884 32652 892
rect 32688 892 32772 912
rect 32688 884 32708 892
rect 32716 884 32744 892
rect 32752 884 32772 892
rect 32808 892 32892 912
rect 32808 884 32828 892
rect 32836 884 32864 892
rect 32872 884 32892 892
rect 32928 892 33012 912
rect 32928 884 32948 892
rect 32956 884 32984 892
rect 32992 884 33012 892
rect 33048 892 33132 912
rect 33048 884 33068 892
rect 33076 884 33104 892
rect 33112 884 33132 892
rect 33168 892 33252 912
rect 33168 884 33188 892
rect 33196 884 33224 892
rect 33232 884 33252 892
rect 33288 892 33372 912
rect 33288 884 33308 892
rect 33316 884 33344 892
rect 33352 884 33372 892
rect 33408 892 33492 912
rect 33408 884 33428 892
rect 33436 884 33464 892
rect 33472 884 33492 892
rect 33528 892 33612 912
rect 33528 884 33548 892
rect 33556 884 33584 892
rect 33592 884 33612 892
rect 33648 892 33732 912
rect 33648 884 33668 892
rect 33676 884 33704 892
rect 33712 884 33732 892
rect 33768 892 33852 912
rect 33768 884 33788 892
rect 33796 884 33824 892
rect 33832 884 33852 892
rect 33888 892 33972 912
rect 33888 884 33908 892
rect 33916 884 33944 892
rect 33952 884 33972 892
rect 34008 892 34092 912
rect 34008 884 34028 892
rect 34036 884 34064 892
rect 34072 884 34092 892
rect 34128 892 34212 912
rect 34128 884 34148 892
rect 34156 884 34184 892
rect 34192 884 34212 892
rect 34248 892 34332 912
rect 34248 884 34268 892
rect 34276 884 34304 892
rect 34312 884 34332 892
rect 34368 892 34452 912
rect 34368 884 34388 892
rect 34396 884 34424 892
rect 34432 884 34452 892
rect 34488 892 34572 912
rect 34488 884 34508 892
rect 34516 884 34544 892
rect 34552 884 34572 892
rect 34608 892 34692 912
rect 34608 884 34628 892
rect 34636 884 34664 892
rect 34672 884 34692 892
rect 34728 892 34812 912
rect 34728 884 34748 892
rect 34756 884 34784 892
rect 34792 884 34812 892
rect 34848 892 34932 912
rect 34848 884 34868 892
rect 34876 884 34904 892
rect 34912 884 34932 892
rect 34968 892 35052 912
rect 34968 884 34988 892
rect 34996 884 35024 892
rect 35032 884 35052 892
rect 35088 892 35172 912
rect 35088 884 35108 892
rect 35116 884 35144 892
rect 35152 884 35172 892
rect 35208 892 35292 912
rect 35208 884 35228 892
rect 35236 884 35264 892
rect 35272 884 35292 892
rect 35328 892 35412 912
rect 35328 884 35348 892
rect 35356 884 35384 892
rect 35392 884 35412 892
rect 35448 892 35532 912
rect 35448 884 35468 892
rect 35476 884 35504 892
rect 35512 884 35532 892
rect 35568 892 35652 912
rect 35568 884 35588 892
rect 35596 884 35624 892
rect 35632 884 35652 892
rect 35688 892 35772 912
rect 35688 884 35708 892
rect 35716 884 35744 892
rect 35752 884 35772 892
rect 35808 892 35892 912
rect 35808 884 35828 892
rect 35836 884 35864 892
rect 35872 884 35892 892
rect 35928 892 36012 912
rect 35928 884 35948 892
rect 35956 884 35984 892
rect 35992 884 36012 892
rect 36048 892 36132 912
rect 36048 884 36068 892
rect 36076 884 36104 892
rect 36112 884 36132 892
rect 36168 892 36252 912
rect 36168 884 36188 892
rect 36196 884 36224 892
rect 36232 884 36252 892
rect 36288 892 36372 912
rect 36288 884 36308 892
rect 36316 884 36344 892
rect 36352 884 36372 892
rect 36408 892 36492 912
rect 36408 884 36428 892
rect 36436 884 36464 892
rect 36472 884 36492 892
rect 36528 892 36612 912
rect 36528 884 36548 892
rect 36556 884 36584 892
rect 36592 884 36612 892
rect 36648 892 36732 912
rect 36648 884 36668 892
rect 36676 884 36704 892
rect 36712 884 36732 892
rect 36768 892 36852 912
rect 36768 884 36788 892
rect 36796 884 36824 892
rect 36832 884 36852 892
rect 36888 892 36972 912
rect 36888 884 36908 892
rect 36916 884 36944 892
rect 36952 884 36972 892
rect 37008 892 37092 912
rect 37008 884 37028 892
rect 37036 884 37064 892
rect 37072 884 37092 892
rect 37128 892 37212 912
rect 37128 884 37148 892
rect 37156 884 37184 892
rect 37192 884 37212 892
rect 37248 892 37332 912
rect 37248 884 37268 892
rect 37276 884 37304 892
rect 37312 884 37332 892
rect 37368 892 37452 912
rect 37368 884 37388 892
rect 37396 884 37424 892
rect 37432 884 37452 892
rect 37488 892 37572 912
rect 37488 884 37508 892
rect 37516 884 37544 892
rect 37552 884 37572 892
rect 37608 892 37692 912
rect 37608 884 37628 892
rect 37636 884 37664 892
rect 37672 884 37692 892
rect 37728 892 37812 912
rect 37728 884 37748 892
rect 37756 884 37784 892
rect 37792 884 37812 892
rect 37848 892 37932 912
rect 37848 884 37868 892
rect 37876 884 37904 892
rect 37912 884 37932 892
rect 37968 892 38052 912
rect 37968 884 37988 892
rect 37996 884 38024 892
rect 38032 884 38052 892
rect 38088 892 38172 912
rect 38088 884 38108 892
rect 38116 884 38144 892
rect 38152 884 38172 892
rect 38208 892 38292 912
rect 38208 884 38228 892
rect 38236 884 38264 892
rect 38272 884 38292 892
rect 38328 892 38412 912
rect 38328 884 38348 892
rect 38356 884 38384 892
rect 38392 884 38412 892
rect 38448 892 38532 912
rect 38448 884 38468 892
rect 38476 884 38504 892
rect 38512 884 38532 892
rect 38568 892 38652 912
rect 38568 884 38588 892
rect 38596 884 38624 892
rect 38632 884 38652 892
rect 38688 892 38772 912
rect 38688 884 38708 892
rect 38716 884 38744 892
rect 38752 884 38772 892
rect 38808 892 38892 912
rect 38808 884 38828 892
rect 38836 884 38864 892
rect 38872 884 38892 892
rect 38928 892 39012 912
rect 38928 884 38948 892
rect 38956 884 38984 892
rect 38992 884 39012 892
rect 39048 892 39132 912
rect 39048 884 39068 892
rect 39076 884 39104 892
rect 39112 884 39132 892
rect 39168 892 39252 912
rect 39168 884 39188 892
rect 39196 884 39224 892
rect 39232 884 39252 892
rect 39288 892 39372 912
rect 39288 884 39308 892
rect 39316 884 39344 892
rect 39352 884 39372 892
rect 39408 892 39492 912
rect 39408 884 39428 892
rect 39436 884 39464 892
rect 39472 884 39492 892
rect 39528 892 39612 912
rect 39528 884 39548 892
rect 39556 884 39584 892
rect 39592 884 39612 892
rect 39648 892 39732 912
rect 39648 884 39668 892
rect 39676 884 39704 892
rect 39712 884 39732 892
rect 39768 892 39852 912
rect 39768 884 39788 892
rect 39796 884 39824 892
rect 39832 884 39852 892
rect 39888 892 39972 912
rect 39888 884 39908 892
rect 39916 884 39944 892
rect 39952 884 39972 892
rect 40008 892 40092 912
rect 40008 884 40028 892
rect 40036 884 40064 892
rect 40072 884 40092 892
rect 40128 892 40212 912
rect 40128 884 40148 892
rect 40156 884 40184 892
rect 40192 884 40212 892
rect 40248 892 40332 912
rect 40248 884 40268 892
rect 40276 884 40304 892
rect 40312 884 40332 892
rect 40368 892 40452 912
rect 40368 884 40388 892
rect 40396 884 40424 892
rect 40432 884 40452 892
rect 40488 892 40572 912
rect 40488 884 40508 892
rect 40516 884 40544 892
rect 40552 884 40572 892
rect 40608 892 40692 912
rect 40608 884 40628 892
rect 40636 884 40664 892
rect 40672 884 40692 892
rect 40728 892 40812 912
rect 40728 884 40748 892
rect 40756 884 40784 892
rect 40792 884 40812 892
rect 40848 892 40932 912
rect 40848 884 40868 892
rect 40876 884 40904 892
rect 40912 884 40932 892
rect 40968 892 41052 912
rect 40968 884 40988 892
rect 40996 884 41024 892
rect 41032 884 41052 892
rect 41088 892 41172 912
rect 41088 884 41108 892
rect 41116 884 41144 892
rect 41152 884 41172 892
rect 41208 892 41292 912
rect 41208 884 41228 892
rect 41236 884 41264 892
rect 41272 884 41292 892
rect 41328 892 41412 912
rect 41328 884 41348 892
rect 41356 884 41384 892
rect 41392 884 41412 892
rect 41448 892 41532 912
rect 41448 884 41468 892
rect 41476 884 41504 892
rect 41512 884 41532 892
rect 41568 892 41652 912
rect 41568 884 41588 892
rect 41596 884 41624 892
rect 41632 884 41652 892
rect 41688 892 41772 912
rect 41688 884 41708 892
rect 41716 884 41744 892
rect 41752 884 41772 892
rect 41808 892 41892 912
rect 41808 884 41828 892
rect 41836 884 41864 892
rect 41872 884 41892 892
rect 41928 892 42012 912
rect 41928 884 41948 892
rect 41956 884 41984 892
rect 41992 884 42012 892
rect 42048 892 42132 912
rect 42048 884 42068 892
rect 42076 884 42104 892
rect 42112 884 42132 892
rect 42168 892 42252 912
rect 42168 884 42188 892
rect 42196 884 42224 892
rect 42232 884 42252 892
rect 42288 892 42372 912
rect 42288 884 42308 892
rect 42316 884 42344 892
rect 42352 884 42372 892
rect 42408 892 42492 912
rect 42408 884 42428 892
rect 42436 884 42464 892
rect 42472 884 42492 892
rect 42528 892 42612 912
rect 42528 884 42548 892
rect 42556 884 42584 892
rect 42592 884 42612 892
rect 42648 892 42732 912
rect 42648 884 42668 892
rect 42676 884 42704 892
rect 42712 884 42732 892
rect 42768 892 42852 912
rect 42768 884 42788 892
rect 42796 884 42824 892
rect 42832 884 42852 892
rect 42888 892 42972 912
rect 42888 884 42908 892
rect 42916 884 42944 892
rect 42952 884 42972 892
rect 43008 892 43092 912
rect 43008 884 43028 892
rect 43036 884 43064 892
rect 43072 884 43092 892
rect 43128 892 43212 912
rect 43128 884 43148 892
rect 43156 884 43184 892
rect 43192 884 43212 892
rect 43248 892 43332 912
rect 43248 884 43268 892
rect 43276 884 43304 892
rect 43312 884 43332 892
rect 43368 892 43452 912
rect 43368 884 43388 892
rect 43396 884 43424 892
rect 43432 884 43452 892
rect 43488 892 43572 912
rect 43488 884 43508 892
rect 43516 884 43544 892
rect 43552 884 43572 892
rect 43608 892 43692 912
rect 43608 884 43628 892
rect 43636 884 43664 892
rect 43672 884 43692 892
rect 43728 892 43812 912
rect 43728 884 43748 892
rect 43756 884 43784 892
rect 43792 884 43812 892
rect 43848 892 43932 912
rect 43848 884 43868 892
rect 43876 884 43904 892
rect 43912 884 43932 892
rect 43968 892 44052 912
rect 43968 884 43988 892
rect 43996 884 44024 892
rect 44032 884 44052 892
rect 44088 892 44172 912
rect 44088 884 44108 892
rect 44116 884 44144 892
rect 44152 884 44172 892
rect 44208 892 44292 912
rect 44208 884 44228 892
rect 44236 884 44264 892
rect 44272 884 44292 892
rect 44328 892 44412 912
rect 44328 884 44348 892
rect 44356 884 44384 892
rect 44392 884 44412 892
rect 44448 892 44532 912
rect 44448 884 44468 892
rect 44476 884 44504 892
rect 44512 884 44532 892
rect 44568 892 44652 912
rect 44568 884 44588 892
rect 44596 884 44624 892
rect 44632 884 44652 892
rect 44688 892 44772 912
rect 44688 884 44708 892
rect 44716 884 44744 892
rect 44752 884 44772 892
rect 44808 892 44892 912
rect 44808 884 44828 892
rect 44836 884 44864 892
rect 44872 884 44892 892
rect 44928 892 45012 912
rect 44928 884 44948 892
rect 44956 884 44984 892
rect 44992 884 45012 892
rect 45048 892 45132 912
rect 45048 884 45068 892
rect 45076 884 45104 892
rect 45112 884 45132 892
rect 45168 892 45252 912
rect 45168 884 45188 892
rect 45196 884 45224 892
rect 45232 884 45252 892
rect 45288 892 45372 912
rect 45288 884 45308 892
rect 45316 884 45344 892
rect 45352 884 45372 892
rect 45408 892 45492 912
rect 45408 884 45428 892
rect 45436 884 45464 892
rect 45472 884 45492 892
rect 45528 892 45612 912
rect 45528 884 45548 892
rect 45556 884 45584 892
rect 45592 884 45612 892
rect 25876 856 25932 884
rect 25996 856 26052 884
rect 26116 856 26172 884
rect 26236 856 26292 884
rect 26356 856 26412 884
rect 26476 856 26532 884
rect 26596 856 26652 884
rect 26716 856 26772 884
rect 26836 856 26892 884
rect 26956 856 27012 884
rect 27076 856 27132 884
rect 27196 856 27252 884
rect 27316 856 27372 884
rect 27436 856 27492 884
rect 27556 856 27612 884
rect 27676 856 27732 884
rect 27796 856 27852 884
rect 27916 856 27972 884
rect 28036 856 28092 884
rect 28156 856 28212 884
rect 28276 856 28332 884
rect 28396 856 28452 884
rect 28516 856 28572 884
rect 28636 856 28692 884
rect 28756 856 28812 884
rect 28876 856 28932 884
rect 28996 856 29052 884
rect 29116 856 29172 884
rect 29236 856 29292 884
rect 29356 856 29412 884
rect 29476 856 29532 884
rect 29596 856 29652 884
rect 29716 856 29772 884
rect 29836 856 29892 884
rect 29956 856 30012 884
rect 30076 856 30132 884
rect 30196 856 30252 884
rect 30316 856 30372 884
rect 30436 856 30492 884
rect 30556 856 30612 884
rect 30676 856 30732 884
rect 30796 856 30852 884
rect 30916 856 30972 884
rect 31036 856 31092 884
rect 31156 856 31212 884
rect 31276 856 31332 884
rect 31396 856 31452 884
rect 31516 856 31572 884
rect 31636 856 31692 884
rect 31756 856 31812 884
rect 31876 856 31932 884
rect 31996 856 32052 884
rect 32116 856 32172 884
rect 32236 856 32292 884
rect 32356 856 32412 884
rect 32476 856 32532 884
rect 32596 856 32652 884
rect 32716 856 32772 884
rect 32836 856 32892 884
rect 32956 856 33012 884
rect 33076 856 33132 884
rect 33196 856 33252 884
rect 33316 856 33372 884
rect 33436 856 33492 884
rect 33556 856 33612 884
rect 33676 856 33732 884
rect 33796 856 33852 884
rect 33916 856 33972 884
rect 34036 856 34092 884
rect 34156 856 34212 884
rect 34276 856 34332 884
rect 34396 856 34452 884
rect 34516 856 34572 884
rect 34636 856 34692 884
rect 34756 856 34812 884
rect 34876 856 34932 884
rect 34996 856 35052 884
rect 35116 856 35172 884
rect 35236 856 35292 884
rect 35356 856 35412 884
rect 35476 856 35532 884
rect 35596 856 35652 884
rect 35716 856 35772 884
rect 35836 856 35892 884
rect 35956 856 36012 884
rect 36076 856 36132 884
rect 36196 856 36252 884
rect 36316 856 36372 884
rect 36436 856 36492 884
rect 36556 856 36612 884
rect 36676 856 36732 884
rect 36796 856 36852 884
rect 36916 856 36972 884
rect 37036 856 37092 884
rect 37156 856 37212 884
rect 37276 856 37332 884
rect 37396 856 37452 884
rect 37516 856 37572 884
rect 37636 856 37692 884
rect 37756 856 37812 884
rect 37876 856 37932 884
rect 37996 856 38052 884
rect 38116 856 38172 884
rect 38236 856 38292 884
rect 38356 856 38412 884
rect 38476 856 38532 884
rect 38596 856 38652 884
rect 38716 856 38772 884
rect 38836 856 38892 884
rect 38956 856 39012 884
rect 39076 856 39132 884
rect 39196 856 39252 884
rect 39316 856 39372 884
rect 39436 856 39492 884
rect 39556 856 39612 884
rect 39676 856 39732 884
rect 39796 856 39852 884
rect 39916 856 39972 884
rect 40036 856 40092 884
rect 40156 856 40212 884
rect 40276 856 40332 884
rect 40396 856 40452 884
rect 40516 856 40572 884
rect 40636 856 40692 884
rect 40756 856 40812 884
rect 40876 856 40932 884
rect 40996 856 41052 884
rect 41116 856 41172 884
rect 41236 856 41292 884
rect 41356 856 41412 884
rect 41476 856 41532 884
rect 41596 856 41652 884
rect 41716 856 41772 884
rect 41836 856 41892 884
rect 41956 856 42012 884
rect 42076 856 42132 884
rect 42196 856 42252 884
rect 42316 856 42372 884
rect 42436 856 42492 884
rect 42556 856 42612 884
rect 42676 856 42732 884
rect 42796 856 42852 884
rect 42916 856 42972 884
rect 43036 856 43092 884
rect 43156 856 43212 884
rect 43276 856 43332 884
rect 43396 856 43452 884
rect 43516 856 43572 884
rect 43636 856 43692 884
rect 43756 856 43812 884
rect 43876 856 43932 884
rect 43996 856 44052 884
rect 44116 856 44172 884
rect 44236 856 44292 884
rect 44356 856 44412 884
rect 44476 856 44532 884
rect 44596 856 44652 884
rect 44716 856 44772 884
rect 44836 856 44892 884
rect 44956 856 45012 884
rect 45076 856 45132 884
rect 45196 856 45252 884
rect 45316 856 45372 884
rect 45436 856 45492 884
rect 45556 856 45612 884
rect 25848 712 25932 732
rect 25848 704 25868 712
rect 25876 704 25904 712
rect 25912 704 25932 712
rect 25968 712 26052 732
rect 25968 704 25988 712
rect 25996 704 26024 712
rect 26032 704 26052 712
rect 26088 712 26172 732
rect 26088 704 26108 712
rect 26116 704 26144 712
rect 26152 704 26172 712
rect 26208 712 26292 732
rect 26208 704 26228 712
rect 26236 704 26264 712
rect 26272 704 26292 712
rect 26328 712 26412 732
rect 26328 704 26348 712
rect 26356 704 26384 712
rect 26392 704 26412 712
rect 26448 712 26532 732
rect 26448 704 26468 712
rect 26476 704 26504 712
rect 26512 704 26532 712
rect 26568 712 26652 732
rect 26568 704 26588 712
rect 26596 704 26624 712
rect 26632 704 26652 712
rect 26688 712 26772 732
rect 26688 704 26708 712
rect 26716 704 26744 712
rect 26752 704 26772 712
rect 26808 712 26892 732
rect 26808 704 26828 712
rect 26836 704 26864 712
rect 26872 704 26892 712
rect 26928 712 27012 732
rect 26928 704 26948 712
rect 26956 704 26984 712
rect 26992 704 27012 712
rect 27048 712 27132 732
rect 27048 704 27068 712
rect 27076 704 27104 712
rect 27112 704 27132 712
rect 27168 712 27252 732
rect 27168 704 27188 712
rect 27196 704 27224 712
rect 27232 704 27252 712
rect 27288 712 27372 732
rect 27288 704 27308 712
rect 27316 704 27344 712
rect 27352 704 27372 712
rect 27408 712 27492 732
rect 27408 704 27428 712
rect 27436 704 27464 712
rect 27472 704 27492 712
rect 27528 712 27612 732
rect 27528 704 27548 712
rect 27556 704 27584 712
rect 27592 704 27612 712
rect 27648 712 27732 732
rect 27648 704 27668 712
rect 27676 704 27704 712
rect 27712 704 27732 712
rect 27768 712 27852 732
rect 27768 704 27788 712
rect 27796 704 27824 712
rect 27832 704 27852 712
rect 27888 712 27972 732
rect 27888 704 27908 712
rect 27916 704 27944 712
rect 27952 704 27972 712
rect 28008 712 28092 732
rect 28008 704 28028 712
rect 28036 704 28064 712
rect 28072 704 28092 712
rect 28128 712 28212 732
rect 28128 704 28148 712
rect 28156 704 28184 712
rect 28192 704 28212 712
rect 28248 712 28332 732
rect 28248 704 28268 712
rect 28276 704 28304 712
rect 28312 704 28332 712
rect 28368 712 28452 732
rect 28368 704 28388 712
rect 28396 704 28424 712
rect 28432 704 28452 712
rect 28488 712 28572 732
rect 28488 704 28508 712
rect 28516 704 28544 712
rect 28552 704 28572 712
rect 28608 712 28692 732
rect 28608 704 28628 712
rect 28636 704 28664 712
rect 28672 704 28692 712
rect 28728 712 28812 732
rect 28728 704 28748 712
rect 28756 704 28784 712
rect 28792 704 28812 712
rect 28848 712 28932 732
rect 28848 704 28868 712
rect 28876 704 28904 712
rect 28912 704 28932 712
rect 28968 712 29052 732
rect 28968 704 28988 712
rect 28996 704 29024 712
rect 29032 704 29052 712
rect 29088 712 29172 732
rect 29088 704 29108 712
rect 29116 704 29144 712
rect 29152 704 29172 712
rect 29208 712 29292 732
rect 29208 704 29228 712
rect 29236 704 29264 712
rect 29272 704 29292 712
rect 29328 712 29412 732
rect 29328 704 29348 712
rect 29356 704 29384 712
rect 29392 704 29412 712
rect 29448 712 29532 732
rect 29448 704 29468 712
rect 29476 704 29504 712
rect 29512 704 29532 712
rect 29568 712 29652 732
rect 29568 704 29588 712
rect 29596 704 29624 712
rect 29632 704 29652 712
rect 29688 712 29772 732
rect 29688 704 29708 712
rect 29716 704 29744 712
rect 29752 704 29772 712
rect 29808 712 29892 732
rect 29808 704 29828 712
rect 29836 704 29864 712
rect 29872 704 29892 712
rect 29928 712 30012 732
rect 29928 704 29948 712
rect 29956 704 29984 712
rect 29992 704 30012 712
rect 30048 712 30132 732
rect 30048 704 30068 712
rect 30076 704 30104 712
rect 30112 704 30132 712
rect 30168 712 30252 732
rect 30168 704 30188 712
rect 30196 704 30224 712
rect 30232 704 30252 712
rect 30288 712 30372 732
rect 30288 704 30308 712
rect 30316 704 30344 712
rect 30352 704 30372 712
rect 30408 712 30492 732
rect 30408 704 30428 712
rect 30436 704 30464 712
rect 30472 704 30492 712
rect 30528 712 30612 732
rect 30528 704 30548 712
rect 30556 704 30584 712
rect 30592 704 30612 712
rect 30648 712 30732 732
rect 30648 704 30668 712
rect 30676 704 30704 712
rect 30712 704 30732 712
rect 30768 712 30852 732
rect 30768 704 30788 712
rect 30796 704 30824 712
rect 30832 704 30852 712
rect 30888 712 30972 732
rect 30888 704 30908 712
rect 30916 704 30944 712
rect 30952 704 30972 712
rect 31008 712 31092 732
rect 31008 704 31028 712
rect 31036 704 31064 712
rect 31072 704 31092 712
rect 31128 712 31212 732
rect 31128 704 31148 712
rect 31156 704 31184 712
rect 31192 704 31212 712
rect 31248 712 31332 732
rect 31248 704 31268 712
rect 31276 704 31304 712
rect 31312 704 31332 712
rect 31368 712 31452 732
rect 31368 704 31388 712
rect 31396 704 31424 712
rect 31432 704 31452 712
rect 31488 712 31572 732
rect 31488 704 31508 712
rect 31516 704 31544 712
rect 31552 704 31572 712
rect 31608 712 31692 732
rect 31608 704 31628 712
rect 31636 704 31664 712
rect 31672 704 31692 712
rect 31728 712 31812 732
rect 31728 704 31748 712
rect 31756 704 31784 712
rect 31792 704 31812 712
rect 31848 712 31932 732
rect 31848 704 31868 712
rect 31876 704 31904 712
rect 31912 704 31932 712
rect 31968 712 32052 732
rect 31968 704 31988 712
rect 31996 704 32024 712
rect 32032 704 32052 712
rect 32088 712 32172 732
rect 32088 704 32108 712
rect 32116 704 32144 712
rect 32152 704 32172 712
rect 32208 712 32292 732
rect 32208 704 32228 712
rect 32236 704 32264 712
rect 32272 704 32292 712
rect 32328 712 32412 732
rect 32328 704 32348 712
rect 32356 704 32384 712
rect 32392 704 32412 712
rect 32448 712 32532 732
rect 32448 704 32468 712
rect 32476 704 32504 712
rect 32512 704 32532 712
rect 32568 712 32652 732
rect 32568 704 32588 712
rect 32596 704 32624 712
rect 32632 704 32652 712
rect 32688 712 32772 732
rect 32688 704 32708 712
rect 32716 704 32744 712
rect 32752 704 32772 712
rect 32808 712 32892 732
rect 32808 704 32828 712
rect 32836 704 32864 712
rect 32872 704 32892 712
rect 32928 712 33012 732
rect 32928 704 32948 712
rect 32956 704 32984 712
rect 32992 704 33012 712
rect 33048 712 33132 732
rect 33048 704 33068 712
rect 33076 704 33104 712
rect 33112 704 33132 712
rect 33168 712 33252 732
rect 33168 704 33188 712
rect 33196 704 33224 712
rect 33232 704 33252 712
rect 33288 712 33372 732
rect 33288 704 33308 712
rect 33316 704 33344 712
rect 33352 704 33372 712
rect 33408 712 33492 732
rect 33408 704 33428 712
rect 33436 704 33464 712
rect 33472 704 33492 712
rect 33528 712 33612 732
rect 33528 704 33548 712
rect 33556 704 33584 712
rect 33592 704 33612 712
rect 33648 712 33732 732
rect 33648 704 33668 712
rect 33676 704 33704 712
rect 33712 704 33732 712
rect 33768 712 33852 732
rect 33768 704 33788 712
rect 33796 704 33824 712
rect 33832 704 33852 712
rect 33888 712 33972 732
rect 33888 704 33908 712
rect 33916 704 33944 712
rect 33952 704 33972 712
rect 34008 712 34092 732
rect 34008 704 34028 712
rect 34036 704 34064 712
rect 34072 704 34092 712
rect 34128 712 34212 732
rect 34128 704 34148 712
rect 34156 704 34184 712
rect 34192 704 34212 712
rect 34248 712 34332 732
rect 34248 704 34268 712
rect 34276 704 34304 712
rect 34312 704 34332 712
rect 34368 712 34452 732
rect 34368 704 34388 712
rect 34396 704 34424 712
rect 34432 704 34452 712
rect 34488 712 34572 732
rect 34488 704 34508 712
rect 34516 704 34544 712
rect 34552 704 34572 712
rect 34608 712 34692 732
rect 34608 704 34628 712
rect 34636 704 34664 712
rect 34672 704 34692 712
rect 34728 712 34812 732
rect 34728 704 34748 712
rect 34756 704 34784 712
rect 34792 704 34812 712
rect 34848 712 34932 732
rect 34848 704 34868 712
rect 34876 704 34904 712
rect 34912 704 34932 712
rect 34968 712 35052 732
rect 34968 704 34988 712
rect 34996 704 35024 712
rect 35032 704 35052 712
rect 35088 712 35172 732
rect 35088 704 35108 712
rect 35116 704 35144 712
rect 35152 704 35172 712
rect 35208 712 35292 732
rect 35208 704 35228 712
rect 35236 704 35264 712
rect 35272 704 35292 712
rect 35328 712 35412 732
rect 35328 704 35348 712
rect 35356 704 35384 712
rect 35392 704 35412 712
rect 35448 712 35532 732
rect 35448 704 35468 712
rect 35476 704 35504 712
rect 35512 704 35532 712
rect 35568 712 35652 732
rect 35568 704 35588 712
rect 35596 704 35624 712
rect 35632 704 35652 712
rect 35688 712 35772 732
rect 35688 704 35708 712
rect 35716 704 35744 712
rect 35752 704 35772 712
rect 35808 712 35892 732
rect 35808 704 35828 712
rect 35836 704 35864 712
rect 35872 704 35892 712
rect 35928 712 36012 732
rect 35928 704 35948 712
rect 35956 704 35984 712
rect 35992 704 36012 712
rect 36048 712 36132 732
rect 36048 704 36068 712
rect 36076 704 36104 712
rect 36112 704 36132 712
rect 36168 712 36252 732
rect 36168 704 36188 712
rect 36196 704 36224 712
rect 36232 704 36252 712
rect 36288 712 36372 732
rect 36288 704 36308 712
rect 36316 704 36344 712
rect 36352 704 36372 712
rect 36408 712 36492 732
rect 36408 704 36428 712
rect 36436 704 36464 712
rect 36472 704 36492 712
rect 36528 712 36612 732
rect 36528 704 36548 712
rect 36556 704 36584 712
rect 36592 704 36612 712
rect 36648 712 36732 732
rect 36648 704 36668 712
rect 36676 704 36704 712
rect 36712 704 36732 712
rect 36768 712 36852 732
rect 36768 704 36788 712
rect 36796 704 36824 712
rect 36832 704 36852 712
rect 36888 712 36972 732
rect 36888 704 36908 712
rect 36916 704 36944 712
rect 36952 704 36972 712
rect 37008 712 37092 732
rect 37008 704 37028 712
rect 37036 704 37064 712
rect 37072 704 37092 712
rect 37128 712 37212 732
rect 37128 704 37148 712
rect 37156 704 37184 712
rect 37192 704 37212 712
rect 37248 712 37332 732
rect 37248 704 37268 712
rect 37276 704 37304 712
rect 37312 704 37332 712
rect 37368 712 37452 732
rect 37368 704 37388 712
rect 37396 704 37424 712
rect 37432 704 37452 712
rect 37488 712 37572 732
rect 37488 704 37508 712
rect 37516 704 37544 712
rect 37552 704 37572 712
rect 37608 712 37692 732
rect 37608 704 37628 712
rect 37636 704 37664 712
rect 37672 704 37692 712
rect 37728 712 37812 732
rect 37728 704 37748 712
rect 37756 704 37784 712
rect 37792 704 37812 712
rect 37848 712 37932 732
rect 37848 704 37868 712
rect 37876 704 37904 712
rect 37912 704 37932 712
rect 37968 712 38052 732
rect 37968 704 37988 712
rect 37996 704 38024 712
rect 38032 704 38052 712
rect 38088 712 38172 732
rect 38088 704 38108 712
rect 38116 704 38144 712
rect 38152 704 38172 712
rect 38208 712 38292 732
rect 38208 704 38228 712
rect 38236 704 38264 712
rect 38272 704 38292 712
rect 38328 712 38412 732
rect 38328 704 38348 712
rect 38356 704 38384 712
rect 38392 704 38412 712
rect 38448 712 38532 732
rect 38448 704 38468 712
rect 38476 704 38504 712
rect 38512 704 38532 712
rect 38568 712 38652 732
rect 38568 704 38588 712
rect 38596 704 38624 712
rect 38632 704 38652 712
rect 38688 712 38772 732
rect 38688 704 38708 712
rect 38716 704 38744 712
rect 38752 704 38772 712
rect 38808 712 38892 732
rect 38808 704 38828 712
rect 38836 704 38864 712
rect 38872 704 38892 712
rect 38928 712 39012 732
rect 38928 704 38948 712
rect 38956 704 38984 712
rect 38992 704 39012 712
rect 39048 712 39132 732
rect 39048 704 39068 712
rect 39076 704 39104 712
rect 39112 704 39132 712
rect 39168 712 39252 732
rect 39168 704 39188 712
rect 39196 704 39224 712
rect 39232 704 39252 712
rect 39288 712 39372 732
rect 39288 704 39308 712
rect 39316 704 39344 712
rect 39352 704 39372 712
rect 39408 712 39492 732
rect 39408 704 39428 712
rect 39436 704 39464 712
rect 39472 704 39492 712
rect 39528 712 39612 732
rect 39528 704 39548 712
rect 39556 704 39584 712
rect 39592 704 39612 712
rect 39648 712 39732 732
rect 39648 704 39668 712
rect 39676 704 39704 712
rect 39712 704 39732 712
rect 39768 712 39852 732
rect 39768 704 39788 712
rect 39796 704 39824 712
rect 39832 704 39852 712
rect 39888 712 39972 732
rect 39888 704 39908 712
rect 39916 704 39944 712
rect 39952 704 39972 712
rect 40008 712 40092 732
rect 40008 704 40028 712
rect 40036 704 40064 712
rect 40072 704 40092 712
rect 40128 712 40212 732
rect 40128 704 40148 712
rect 40156 704 40184 712
rect 40192 704 40212 712
rect 40248 712 40332 732
rect 40248 704 40268 712
rect 40276 704 40304 712
rect 40312 704 40332 712
rect 40368 712 40452 732
rect 40368 704 40388 712
rect 40396 704 40424 712
rect 40432 704 40452 712
rect 40488 712 40572 732
rect 40488 704 40508 712
rect 40516 704 40544 712
rect 40552 704 40572 712
rect 40608 712 40692 732
rect 40608 704 40628 712
rect 40636 704 40664 712
rect 40672 704 40692 712
rect 40728 712 40812 732
rect 40728 704 40748 712
rect 40756 704 40784 712
rect 40792 704 40812 712
rect 40848 712 40932 732
rect 40848 704 40868 712
rect 40876 704 40904 712
rect 40912 704 40932 712
rect 40968 712 41052 732
rect 40968 704 40988 712
rect 40996 704 41024 712
rect 41032 704 41052 712
rect 41088 712 41172 732
rect 41088 704 41108 712
rect 41116 704 41144 712
rect 41152 704 41172 712
rect 41208 712 41292 732
rect 41208 704 41228 712
rect 41236 704 41264 712
rect 41272 704 41292 712
rect 41328 712 41412 732
rect 41328 704 41348 712
rect 41356 704 41384 712
rect 41392 704 41412 712
rect 41448 712 41532 732
rect 41448 704 41468 712
rect 41476 704 41504 712
rect 41512 704 41532 712
rect 41568 712 41652 732
rect 41568 704 41588 712
rect 41596 704 41624 712
rect 41632 704 41652 712
rect 41688 712 41772 732
rect 41688 704 41708 712
rect 41716 704 41744 712
rect 41752 704 41772 712
rect 41808 712 41892 732
rect 41808 704 41828 712
rect 41836 704 41864 712
rect 41872 704 41892 712
rect 41928 712 42012 732
rect 41928 704 41948 712
rect 41956 704 41984 712
rect 41992 704 42012 712
rect 42048 712 42132 732
rect 42048 704 42068 712
rect 42076 704 42104 712
rect 42112 704 42132 712
rect 42168 712 42252 732
rect 42168 704 42188 712
rect 42196 704 42224 712
rect 42232 704 42252 712
rect 42288 712 42372 732
rect 42288 704 42308 712
rect 42316 704 42344 712
rect 42352 704 42372 712
rect 42408 712 42492 732
rect 42408 704 42428 712
rect 42436 704 42464 712
rect 42472 704 42492 712
rect 42528 712 42612 732
rect 42528 704 42548 712
rect 42556 704 42584 712
rect 42592 704 42612 712
rect 42648 712 42732 732
rect 42648 704 42668 712
rect 42676 704 42704 712
rect 42712 704 42732 712
rect 42768 712 42852 732
rect 42768 704 42788 712
rect 42796 704 42824 712
rect 42832 704 42852 712
rect 42888 712 42972 732
rect 42888 704 42908 712
rect 42916 704 42944 712
rect 42952 704 42972 712
rect 43008 712 43092 732
rect 43008 704 43028 712
rect 43036 704 43064 712
rect 43072 704 43092 712
rect 43128 712 43212 732
rect 43128 704 43148 712
rect 43156 704 43184 712
rect 43192 704 43212 712
rect 43248 712 43332 732
rect 43248 704 43268 712
rect 43276 704 43304 712
rect 43312 704 43332 712
rect 43368 712 43452 732
rect 43368 704 43388 712
rect 43396 704 43424 712
rect 43432 704 43452 712
rect 43488 712 43572 732
rect 43488 704 43508 712
rect 43516 704 43544 712
rect 43552 704 43572 712
rect 43608 712 43692 732
rect 43608 704 43628 712
rect 43636 704 43664 712
rect 43672 704 43692 712
rect 43728 712 43812 732
rect 43728 704 43748 712
rect 43756 704 43784 712
rect 43792 704 43812 712
rect 43848 712 43932 732
rect 43848 704 43868 712
rect 43876 704 43904 712
rect 43912 704 43932 712
rect 43968 712 44052 732
rect 43968 704 43988 712
rect 43996 704 44024 712
rect 44032 704 44052 712
rect 44088 712 44172 732
rect 44088 704 44108 712
rect 44116 704 44144 712
rect 44152 704 44172 712
rect 44208 712 44292 732
rect 44208 704 44228 712
rect 44236 704 44264 712
rect 44272 704 44292 712
rect 44328 712 44412 732
rect 44328 704 44348 712
rect 44356 704 44384 712
rect 44392 704 44412 712
rect 44448 712 44532 732
rect 44448 704 44468 712
rect 44476 704 44504 712
rect 44512 704 44532 712
rect 44568 712 44652 732
rect 44568 704 44588 712
rect 44596 704 44624 712
rect 44632 704 44652 712
rect 44688 712 44772 732
rect 44688 704 44708 712
rect 44716 704 44744 712
rect 44752 704 44772 712
rect 44808 712 44892 732
rect 44808 704 44828 712
rect 44836 704 44864 712
rect 44872 704 44892 712
rect 44928 712 45012 732
rect 44928 704 44948 712
rect 44956 704 44984 712
rect 44992 704 45012 712
rect 45048 712 45132 732
rect 45048 704 45068 712
rect 45076 704 45104 712
rect 45112 704 45132 712
rect 45168 712 45252 732
rect 45168 704 45188 712
rect 45196 704 45224 712
rect 45232 704 45252 712
rect 45288 712 45372 732
rect 45288 704 45308 712
rect 45316 704 45344 712
rect 45352 704 45372 712
rect 45408 712 45492 732
rect 45408 704 45428 712
rect 45436 704 45464 712
rect 45472 704 45492 712
rect 45528 712 45612 732
rect 45528 704 45548 712
rect 45556 704 45584 712
rect 45592 704 45612 712
rect 25876 676 25932 704
rect 25996 676 26052 704
rect 26116 676 26172 704
rect 26236 676 26292 704
rect 26356 676 26412 704
rect 26476 676 26532 704
rect 26596 676 26652 704
rect 26716 676 26772 704
rect 26836 676 26892 704
rect 26956 676 27012 704
rect 27076 676 27132 704
rect 27196 676 27252 704
rect 27316 676 27372 704
rect 27436 676 27492 704
rect 27556 676 27612 704
rect 27676 676 27732 704
rect 27796 676 27852 704
rect 27916 676 27972 704
rect 28036 676 28092 704
rect 28156 676 28212 704
rect 28276 676 28332 704
rect 28396 676 28452 704
rect 28516 676 28572 704
rect 28636 676 28692 704
rect 28756 676 28812 704
rect 28876 676 28932 704
rect 28996 676 29052 704
rect 29116 676 29172 704
rect 29236 676 29292 704
rect 29356 676 29412 704
rect 29476 676 29532 704
rect 29596 676 29652 704
rect 29716 676 29772 704
rect 29836 676 29892 704
rect 29956 676 30012 704
rect 30076 676 30132 704
rect 30196 676 30252 704
rect 30316 676 30372 704
rect 30436 676 30492 704
rect 30556 676 30612 704
rect 30676 676 30732 704
rect 30796 676 30852 704
rect 30916 676 30972 704
rect 31036 676 31092 704
rect 31156 676 31212 704
rect 31276 676 31332 704
rect 31396 676 31452 704
rect 31516 676 31572 704
rect 31636 676 31692 704
rect 31756 676 31812 704
rect 31876 676 31932 704
rect 31996 676 32052 704
rect 32116 676 32172 704
rect 32236 676 32292 704
rect 32356 676 32412 704
rect 32476 676 32532 704
rect 32596 676 32652 704
rect 32716 676 32772 704
rect 32836 676 32892 704
rect 32956 676 33012 704
rect 33076 676 33132 704
rect 33196 676 33252 704
rect 33316 676 33372 704
rect 33436 676 33492 704
rect 33556 676 33612 704
rect 33676 676 33732 704
rect 33796 676 33852 704
rect 33916 676 33972 704
rect 34036 676 34092 704
rect 34156 676 34212 704
rect 34276 676 34332 704
rect 34396 676 34452 704
rect 34516 676 34572 704
rect 34636 676 34692 704
rect 34756 676 34812 704
rect 34876 676 34932 704
rect 34996 676 35052 704
rect 35116 676 35172 704
rect 35236 676 35292 704
rect 35356 676 35412 704
rect 35476 676 35532 704
rect 35596 676 35652 704
rect 35716 676 35772 704
rect 35836 676 35892 704
rect 35956 676 36012 704
rect 36076 676 36132 704
rect 36196 676 36252 704
rect 36316 676 36372 704
rect 36436 676 36492 704
rect 36556 676 36612 704
rect 36676 676 36732 704
rect 36796 676 36852 704
rect 36916 676 36972 704
rect 37036 676 37092 704
rect 37156 676 37212 704
rect 37276 676 37332 704
rect 37396 676 37452 704
rect 37516 676 37572 704
rect 37636 676 37692 704
rect 37756 676 37812 704
rect 37876 676 37932 704
rect 37996 676 38052 704
rect 38116 676 38172 704
rect 38236 676 38292 704
rect 38356 676 38412 704
rect 38476 676 38532 704
rect 38596 676 38652 704
rect 38716 676 38772 704
rect 38836 676 38892 704
rect 38956 676 39012 704
rect 39076 676 39132 704
rect 39196 676 39252 704
rect 39316 676 39372 704
rect 39436 676 39492 704
rect 39556 676 39612 704
rect 39676 676 39732 704
rect 39796 676 39852 704
rect 39916 676 39972 704
rect 40036 676 40092 704
rect 40156 676 40212 704
rect 40276 676 40332 704
rect 40396 676 40452 704
rect 40516 676 40572 704
rect 40636 676 40692 704
rect 40756 676 40812 704
rect 40876 676 40932 704
rect 40996 676 41052 704
rect 41116 676 41172 704
rect 41236 676 41292 704
rect 41356 676 41412 704
rect 41476 676 41532 704
rect 41596 676 41652 704
rect 41716 676 41772 704
rect 41836 676 41892 704
rect 41956 676 42012 704
rect 42076 676 42132 704
rect 42196 676 42252 704
rect 42316 676 42372 704
rect 42436 676 42492 704
rect 42556 676 42612 704
rect 42676 676 42732 704
rect 42796 676 42852 704
rect 42916 676 42972 704
rect 43036 676 43092 704
rect 43156 676 43212 704
rect 43276 676 43332 704
rect 43396 676 43452 704
rect 43516 676 43572 704
rect 43636 676 43692 704
rect 43756 676 43812 704
rect 43876 676 43932 704
rect 43996 676 44052 704
rect 44116 676 44172 704
rect 44236 676 44292 704
rect 44356 676 44412 704
rect 44476 676 44532 704
rect 44596 676 44652 704
rect 44716 676 44772 704
rect 44836 676 44892 704
rect 44956 676 45012 704
rect 45076 676 45132 704
rect 45196 676 45252 704
rect 45316 676 45372 704
rect 45436 676 45492 704
rect 45556 676 45612 704
rect 25848 532 25932 552
rect 25848 524 25868 532
rect 25876 524 25904 532
rect 25912 524 25932 532
rect 25968 532 26052 552
rect 25968 524 25988 532
rect 25996 524 26024 532
rect 26032 524 26052 532
rect 26088 532 26172 552
rect 26088 524 26108 532
rect 26116 524 26144 532
rect 26152 524 26172 532
rect 26208 532 26292 552
rect 26208 524 26228 532
rect 26236 524 26264 532
rect 26272 524 26292 532
rect 26328 532 26412 552
rect 26328 524 26348 532
rect 26356 524 26384 532
rect 26392 524 26412 532
rect 26448 532 26532 552
rect 26448 524 26468 532
rect 26476 524 26504 532
rect 26512 524 26532 532
rect 26568 532 26652 552
rect 26568 524 26588 532
rect 26596 524 26624 532
rect 26632 524 26652 532
rect 26688 532 26772 552
rect 26688 524 26708 532
rect 26716 524 26744 532
rect 26752 524 26772 532
rect 26808 532 26892 552
rect 26808 524 26828 532
rect 26836 524 26864 532
rect 26872 524 26892 532
rect 26928 532 27012 552
rect 26928 524 26948 532
rect 26956 524 26984 532
rect 26992 524 27012 532
rect 27048 532 27132 552
rect 27048 524 27068 532
rect 27076 524 27104 532
rect 27112 524 27132 532
rect 27168 532 27252 552
rect 27168 524 27188 532
rect 27196 524 27224 532
rect 27232 524 27252 532
rect 27288 532 27372 552
rect 27288 524 27308 532
rect 27316 524 27344 532
rect 27352 524 27372 532
rect 27408 532 27492 552
rect 27408 524 27428 532
rect 27436 524 27464 532
rect 27472 524 27492 532
rect 27528 532 27612 552
rect 27528 524 27548 532
rect 27556 524 27584 532
rect 27592 524 27612 532
rect 27648 532 27732 552
rect 27648 524 27668 532
rect 27676 524 27704 532
rect 27712 524 27732 532
rect 27768 532 27852 552
rect 27768 524 27788 532
rect 27796 524 27824 532
rect 27832 524 27852 532
rect 27888 532 27972 552
rect 27888 524 27908 532
rect 27916 524 27944 532
rect 27952 524 27972 532
rect 28008 532 28092 552
rect 28008 524 28028 532
rect 28036 524 28064 532
rect 28072 524 28092 532
rect 28128 532 28212 552
rect 28128 524 28148 532
rect 28156 524 28184 532
rect 28192 524 28212 532
rect 28248 532 28332 552
rect 28248 524 28268 532
rect 28276 524 28304 532
rect 28312 524 28332 532
rect 28368 532 28452 552
rect 28368 524 28388 532
rect 28396 524 28424 532
rect 28432 524 28452 532
rect 28488 532 28572 552
rect 28488 524 28508 532
rect 28516 524 28544 532
rect 28552 524 28572 532
rect 28608 532 28692 552
rect 28608 524 28628 532
rect 28636 524 28664 532
rect 28672 524 28692 532
rect 28728 532 28812 552
rect 28728 524 28748 532
rect 28756 524 28784 532
rect 28792 524 28812 532
rect 28848 532 28932 552
rect 28848 524 28868 532
rect 28876 524 28904 532
rect 28912 524 28932 532
rect 28968 532 29052 552
rect 28968 524 28988 532
rect 28996 524 29024 532
rect 29032 524 29052 532
rect 29088 532 29172 552
rect 29088 524 29108 532
rect 29116 524 29144 532
rect 29152 524 29172 532
rect 29208 532 29292 552
rect 29208 524 29228 532
rect 29236 524 29264 532
rect 29272 524 29292 532
rect 29328 532 29412 552
rect 29328 524 29348 532
rect 29356 524 29384 532
rect 29392 524 29412 532
rect 29448 532 29532 552
rect 29448 524 29468 532
rect 29476 524 29504 532
rect 29512 524 29532 532
rect 29568 532 29652 552
rect 29568 524 29588 532
rect 29596 524 29624 532
rect 29632 524 29652 532
rect 29688 532 29772 552
rect 29688 524 29708 532
rect 29716 524 29744 532
rect 29752 524 29772 532
rect 29808 532 29892 552
rect 29808 524 29828 532
rect 29836 524 29864 532
rect 29872 524 29892 532
rect 29928 532 30012 552
rect 29928 524 29948 532
rect 29956 524 29984 532
rect 29992 524 30012 532
rect 30048 532 30132 552
rect 30048 524 30068 532
rect 30076 524 30104 532
rect 30112 524 30132 532
rect 30168 532 30252 552
rect 30168 524 30188 532
rect 30196 524 30224 532
rect 30232 524 30252 532
rect 30288 532 30372 552
rect 30288 524 30308 532
rect 30316 524 30344 532
rect 30352 524 30372 532
rect 30408 532 30492 552
rect 30408 524 30428 532
rect 30436 524 30464 532
rect 30472 524 30492 532
rect 30528 532 30612 552
rect 30528 524 30548 532
rect 30556 524 30584 532
rect 30592 524 30612 532
rect 30648 532 30732 552
rect 30648 524 30668 532
rect 30676 524 30704 532
rect 30712 524 30732 532
rect 30768 532 30852 552
rect 30768 524 30788 532
rect 30796 524 30824 532
rect 30832 524 30852 532
rect 30888 532 30972 552
rect 30888 524 30908 532
rect 30916 524 30944 532
rect 30952 524 30972 532
rect 31008 532 31092 552
rect 31008 524 31028 532
rect 31036 524 31064 532
rect 31072 524 31092 532
rect 31128 532 31212 552
rect 31128 524 31148 532
rect 31156 524 31184 532
rect 31192 524 31212 532
rect 31248 532 31332 552
rect 31248 524 31268 532
rect 31276 524 31304 532
rect 31312 524 31332 532
rect 31368 532 31452 552
rect 31368 524 31388 532
rect 31396 524 31424 532
rect 31432 524 31452 532
rect 31488 532 31572 552
rect 31488 524 31508 532
rect 31516 524 31544 532
rect 31552 524 31572 532
rect 31608 532 31692 552
rect 31608 524 31628 532
rect 31636 524 31664 532
rect 31672 524 31692 532
rect 31728 532 31812 552
rect 31728 524 31748 532
rect 31756 524 31784 532
rect 31792 524 31812 532
rect 31848 532 31932 552
rect 31848 524 31868 532
rect 31876 524 31904 532
rect 31912 524 31932 532
rect 31968 532 32052 552
rect 31968 524 31988 532
rect 31996 524 32024 532
rect 32032 524 32052 532
rect 32088 532 32172 552
rect 32088 524 32108 532
rect 32116 524 32144 532
rect 32152 524 32172 532
rect 32208 532 32292 552
rect 32208 524 32228 532
rect 32236 524 32264 532
rect 32272 524 32292 532
rect 32328 532 32412 552
rect 32328 524 32348 532
rect 32356 524 32384 532
rect 32392 524 32412 532
rect 32448 532 32532 552
rect 32448 524 32468 532
rect 32476 524 32504 532
rect 32512 524 32532 532
rect 32568 532 32652 552
rect 32568 524 32588 532
rect 32596 524 32624 532
rect 32632 524 32652 532
rect 32688 532 32772 552
rect 32688 524 32708 532
rect 32716 524 32744 532
rect 32752 524 32772 532
rect 32808 532 32892 552
rect 32808 524 32828 532
rect 32836 524 32864 532
rect 32872 524 32892 532
rect 32928 532 33012 552
rect 32928 524 32948 532
rect 32956 524 32984 532
rect 32992 524 33012 532
rect 33048 532 33132 552
rect 33048 524 33068 532
rect 33076 524 33104 532
rect 33112 524 33132 532
rect 33168 532 33252 552
rect 33168 524 33188 532
rect 33196 524 33224 532
rect 33232 524 33252 532
rect 33288 532 33372 552
rect 33288 524 33308 532
rect 33316 524 33344 532
rect 33352 524 33372 532
rect 33408 532 33492 552
rect 33408 524 33428 532
rect 33436 524 33464 532
rect 33472 524 33492 532
rect 33528 532 33612 552
rect 33528 524 33548 532
rect 33556 524 33584 532
rect 33592 524 33612 532
rect 33648 532 33732 552
rect 33648 524 33668 532
rect 33676 524 33704 532
rect 33712 524 33732 532
rect 33768 532 33852 552
rect 33768 524 33788 532
rect 33796 524 33824 532
rect 33832 524 33852 532
rect 33888 532 33972 552
rect 33888 524 33908 532
rect 33916 524 33944 532
rect 33952 524 33972 532
rect 34008 532 34092 552
rect 34008 524 34028 532
rect 34036 524 34064 532
rect 34072 524 34092 532
rect 34128 532 34212 552
rect 34128 524 34148 532
rect 34156 524 34184 532
rect 34192 524 34212 532
rect 34248 532 34332 552
rect 34248 524 34268 532
rect 34276 524 34304 532
rect 34312 524 34332 532
rect 34368 532 34452 552
rect 34368 524 34388 532
rect 34396 524 34424 532
rect 34432 524 34452 532
rect 34488 532 34572 552
rect 34488 524 34508 532
rect 34516 524 34544 532
rect 34552 524 34572 532
rect 34608 532 34692 552
rect 34608 524 34628 532
rect 34636 524 34664 532
rect 34672 524 34692 532
rect 34728 532 34812 552
rect 34728 524 34748 532
rect 34756 524 34784 532
rect 34792 524 34812 532
rect 34848 532 34932 552
rect 34848 524 34868 532
rect 34876 524 34904 532
rect 34912 524 34932 532
rect 34968 532 35052 552
rect 34968 524 34988 532
rect 34996 524 35024 532
rect 35032 524 35052 532
rect 35088 532 35172 552
rect 35088 524 35108 532
rect 35116 524 35144 532
rect 35152 524 35172 532
rect 35208 532 35292 552
rect 35208 524 35228 532
rect 35236 524 35264 532
rect 35272 524 35292 532
rect 35328 532 35412 552
rect 35328 524 35348 532
rect 35356 524 35384 532
rect 35392 524 35412 532
rect 35448 532 35532 552
rect 35448 524 35468 532
rect 35476 524 35504 532
rect 35512 524 35532 532
rect 35568 532 35652 552
rect 35568 524 35588 532
rect 35596 524 35624 532
rect 35632 524 35652 532
rect 35688 532 35772 552
rect 35688 524 35708 532
rect 35716 524 35744 532
rect 35752 524 35772 532
rect 35808 532 35892 552
rect 35808 524 35828 532
rect 35836 524 35864 532
rect 35872 524 35892 532
rect 35928 532 36012 552
rect 35928 524 35948 532
rect 35956 524 35984 532
rect 35992 524 36012 532
rect 36048 532 36132 552
rect 36048 524 36068 532
rect 36076 524 36104 532
rect 36112 524 36132 532
rect 36168 532 36252 552
rect 36168 524 36188 532
rect 36196 524 36224 532
rect 36232 524 36252 532
rect 36288 532 36372 552
rect 36288 524 36308 532
rect 36316 524 36344 532
rect 36352 524 36372 532
rect 36408 532 36492 552
rect 36408 524 36428 532
rect 36436 524 36464 532
rect 36472 524 36492 532
rect 36528 532 36612 552
rect 36528 524 36548 532
rect 36556 524 36584 532
rect 36592 524 36612 532
rect 36648 532 36732 552
rect 36648 524 36668 532
rect 36676 524 36704 532
rect 36712 524 36732 532
rect 36768 532 36852 552
rect 36768 524 36788 532
rect 36796 524 36824 532
rect 36832 524 36852 532
rect 36888 532 36972 552
rect 36888 524 36908 532
rect 36916 524 36944 532
rect 36952 524 36972 532
rect 37008 532 37092 552
rect 37008 524 37028 532
rect 37036 524 37064 532
rect 37072 524 37092 532
rect 37128 532 37212 552
rect 37128 524 37148 532
rect 37156 524 37184 532
rect 37192 524 37212 532
rect 37248 532 37332 552
rect 37248 524 37268 532
rect 37276 524 37304 532
rect 37312 524 37332 532
rect 37368 532 37452 552
rect 37368 524 37388 532
rect 37396 524 37424 532
rect 37432 524 37452 532
rect 37488 532 37572 552
rect 37488 524 37508 532
rect 37516 524 37544 532
rect 37552 524 37572 532
rect 37608 532 37692 552
rect 37608 524 37628 532
rect 37636 524 37664 532
rect 37672 524 37692 532
rect 37728 532 37812 552
rect 37728 524 37748 532
rect 37756 524 37784 532
rect 37792 524 37812 532
rect 37848 532 37932 552
rect 37848 524 37868 532
rect 37876 524 37904 532
rect 37912 524 37932 532
rect 37968 532 38052 552
rect 37968 524 37988 532
rect 37996 524 38024 532
rect 38032 524 38052 532
rect 38088 532 38172 552
rect 38088 524 38108 532
rect 38116 524 38144 532
rect 38152 524 38172 532
rect 38208 532 38292 552
rect 38208 524 38228 532
rect 38236 524 38264 532
rect 38272 524 38292 532
rect 38328 532 38412 552
rect 38328 524 38348 532
rect 38356 524 38384 532
rect 38392 524 38412 532
rect 38448 532 38532 552
rect 38448 524 38468 532
rect 38476 524 38504 532
rect 38512 524 38532 532
rect 38568 532 38652 552
rect 38568 524 38588 532
rect 38596 524 38624 532
rect 38632 524 38652 532
rect 38688 532 38772 552
rect 38688 524 38708 532
rect 38716 524 38744 532
rect 38752 524 38772 532
rect 38808 532 38892 552
rect 38808 524 38828 532
rect 38836 524 38864 532
rect 38872 524 38892 532
rect 38928 532 39012 552
rect 38928 524 38948 532
rect 38956 524 38984 532
rect 38992 524 39012 532
rect 39048 532 39132 552
rect 39048 524 39068 532
rect 39076 524 39104 532
rect 39112 524 39132 532
rect 39168 532 39252 552
rect 39168 524 39188 532
rect 39196 524 39224 532
rect 39232 524 39252 532
rect 39288 532 39372 552
rect 39288 524 39308 532
rect 39316 524 39344 532
rect 39352 524 39372 532
rect 39408 532 39492 552
rect 39408 524 39428 532
rect 39436 524 39464 532
rect 39472 524 39492 532
rect 39528 532 39612 552
rect 39528 524 39548 532
rect 39556 524 39584 532
rect 39592 524 39612 532
rect 39648 532 39732 552
rect 39648 524 39668 532
rect 39676 524 39704 532
rect 39712 524 39732 532
rect 39768 532 39852 552
rect 39768 524 39788 532
rect 39796 524 39824 532
rect 39832 524 39852 532
rect 39888 532 39972 552
rect 39888 524 39908 532
rect 39916 524 39944 532
rect 39952 524 39972 532
rect 40008 532 40092 552
rect 40008 524 40028 532
rect 40036 524 40064 532
rect 40072 524 40092 532
rect 40128 532 40212 552
rect 40128 524 40148 532
rect 40156 524 40184 532
rect 40192 524 40212 532
rect 40248 532 40332 552
rect 40248 524 40268 532
rect 40276 524 40304 532
rect 40312 524 40332 532
rect 40368 532 40452 552
rect 40368 524 40388 532
rect 40396 524 40424 532
rect 40432 524 40452 532
rect 40488 532 40572 552
rect 40488 524 40508 532
rect 40516 524 40544 532
rect 40552 524 40572 532
rect 40608 532 40692 552
rect 40608 524 40628 532
rect 40636 524 40664 532
rect 40672 524 40692 532
rect 40728 532 40812 552
rect 40728 524 40748 532
rect 40756 524 40784 532
rect 40792 524 40812 532
rect 40848 532 40932 552
rect 40848 524 40868 532
rect 40876 524 40904 532
rect 40912 524 40932 532
rect 40968 532 41052 552
rect 40968 524 40988 532
rect 40996 524 41024 532
rect 41032 524 41052 532
rect 41088 532 41172 552
rect 41088 524 41108 532
rect 41116 524 41144 532
rect 41152 524 41172 532
rect 41208 532 41292 552
rect 41208 524 41228 532
rect 41236 524 41264 532
rect 41272 524 41292 532
rect 41328 532 41412 552
rect 41328 524 41348 532
rect 41356 524 41384 532
rect 41392 524 41412 532
rect 41448 532 41532 552
rect 41448 524 41468 532
rect 41476 524 41504 532
rect 41512 524 41532 532
rect 41568 532 41652 552
rect 41568 524 41588 532
rect 41596 524 41624 532
rect 41632 524 41652 532
rect 41688 532 41772 552
rect 41688 524 41708 532
rect 41716 524 41744 532
rect 41752 524 41772 532
rect 41808 532 41892 552
rect 41808 524 41828 532
rect 41836 524 41864 532
rect 41872 524 41892 532
rect 41928 532 42012 552
rect 41928 524 41948 532
rect 41956 524 41984 532
rect 41992 524 42012 532
rect 42048 532 42132 552
rect 42048 524 42068 532
rect 42076 524 42104 532
rect 42112 524 42132 532
rect 42168 532 42252 552
rect 42168 524 42188 532
rect 42196 524 42224 532
rect 42232 524 42252 532
rect 42288 532 42372 552
rect 42288 524 42308 532
rect 42316 524 42344 532
rect 42352 524 42372 532
rect 42408 532 42492 552
rect 42408 524 42428 532
rect 42436 524 42464 532
rect 42472 524 42492 532
rect 42528 532 42612 552
rect 42528 524 42548 532
rect 42556 524 42584 532
rect 42592 524 42612 532
rect 42648 532 42732 552
rect 42648 524 42668 532
rect 42676 524 42704 532
rect 42712 524 42732 532
rect 42768 532 42852 552
rect 42768 524 42788 532
rect 42796 524 42824 532
rect 42832 524 42852 532
rect 42888 532 42972 552
rect 42888 524 42908 532
rect 42916 524 42944 532
rect 42952 524 42972 532
rect 43008 532 43092 552
rect 43008 524 43028 532
rect 43036 524 43064 532
rect 43072 524 43092 532
rect 43128 532 43212 552
rect 43128 524 43148 532
rect 43156 524 43184 532
rect 43192 524 43212 532
rect 43248 532 43332 552
rect 43248 524 43268 532
rect 43276 524 43304 532
rect 43312 524 43332 532
rect 43368 532 43452 552
rect 43368 524 43388 532
rect 43396 524 43424 532
rect 43432 524 43452 532
rect 43488 532 43572 552
rect 43488 524 43508 532
rect 43516 524 43544 532
rect 43552 524 43572 532
rect 43608 532 43692 552
rect 43608 524 43628 532
rect 43636 524 43664 532
rect 43672 524 43692 532
rect 43728 532 43812 552
rect 43728 524 43748 532
rect 43756 524 43784 532
rect 43792 524 43812 532
rect 43848 532 43932 552
rect 43848 524 43868 532
rect 43876 524 43904 532
rect 43912 524 43932 532
rect 43968 532 44052 552
rect 43968 524 43988 532
rect 43996 524 44024 532
rect 44032 524 44052 532
rect 44088 532 44172 552
rect 44088 524 44108 532
rect 44116 524 44144 532
rect 44152 524 44172 532
rect 44208 532 44292 552
rect 44208 524 44228 532
rect 44236 524 44264 532
rect 44272 524 44292 532
rect 44328 532 44412 552
rect 44328 524 44348 532
rect 44356 524 44384 532
rect 44392 524 44412 532
rect 44448 532 44532 552
rect 44448 524 44468 532
rect 44476 524 44504 532
rect 44512 524 44532 532
rect 44568 532 44652 552
rect 44568 524 44588 532
rect 44596 524 44624 532
rect 44632 524 44652 532
rect 44688 532 44772 552
rect 44688 524 44708 532
rect 44716 524 44744 532
rect 44752 524 44772 532
rect 44808 532 44892 552
rect 44808 524 44828 532
rect 44836 524 44864 532
rect 44872 524 44892 532
rect 44928 532 45012 552
rect 44928 524 44948 532
rect 44956 524 44984 532
rect 44992 524 45012 532
rect 45048 532 45132 552
rect 45048 524 45068 532
rect 45076 524 45104 532
rect 45112 524 45132 532
rect 45168 532 45252 552
rect 45168 524 45188 532
rect 45196 524 45224 532
rect 45232 524 45252 532
rect 45288 532 45372 552
rect 45288 524 45308 532
rect 45316 524 45344 532
rect 45352 524 45372 532
rect 45408 532 45492 552
rect 45408 524 45428 532
rect 45436 524 45464 532
rect 45472 524 45492 532
rect 45528 532 45612 552
rect 45528 524 45548 532
rect 45556 524 45584 532
rect 45592 524 45612 532
rect 25876 496 25932 524
rect 25996 496 26052 524
rect 26116 496 26172 524
rect 26236 496 26292 524
rect 26356 496 26412 524
rect 26476 496 26532 524
rect 26596 496 26652 524
rect 26716 496 26772 524
rect 26836 496 26892 524
rect 26956 496 27012 524
rect 27076 496 27132 524
rect 27196 496 27252 524
rect 27316 496 27372 524
rect 27436 496 27492 524
rect 27556 496 27612 524
rect 27676 496 27732 524
rect 27796 496 27852 524
rect 27916 496 27972 524
rect 28036 496 28092 524
rect 28156 496 28212 524
rect 28276 496 28332 524
rect 28396 496 28452 524
rect 28516 496 28572 524
rect 28636 496 28692 524
rect 28756 496 28812 524
rect 28876 496 28932 524
rect 28996 496 29052 524
rect 29116 496 29172 524
rect 29236 496 29292 524
rect 29356 496 29412 524
rect 29476 496 29532 524
rect 29596 496 29652 524
rect 29716 496 29772 524
rect 29836 496 29892 524
rect 29956 496 30012 524
rect 30076 496 30132 524
rect 30196 496 30252 524
rect 30316 496 30372 524
rect 30436 496 30492 524
rect 30556 496 30612 524
rect 30676 496 30732 524
rect 30796 496 30852 524
rect 30916 496 30972 524
rect 31036 496 31092 524
rect 31156 496 31212 524
rect 31276 496 31332 524
rect 31396 496 31452 524
rect 31516 496 31572 524
rect 31636 496 31692 524
rect 31756 496 31812 524
rect 31876 496 31932 524
rect 31996 496 32052 524
rect 32116 496 32172 524
rect 32236 496 32292 524
rect 32356 496 32412 524
rect 32476 496 32532 524
rect 32596 496 32652 524
rect 32716 496 32772 524
rect 32836 496 32892 524
rect 32956 496 33012 524
rect 33076 496 33132 524
rect 33196 496 33252 524
rect 33316 496 33372 524
rect 33436 496 33492 524
rect 33556 496 33612 524
rect 33676 496 33732 524
rect 33796 496 33852 524
rect 33916 496 33972 524
rect 34036 496 34092 524
rect 34156 496 34212 524
rect 34276 496 34332 524
rect 34396 496 34452 524
rect 34516 496 34572 524
rect 34636 496 34692 524
rect 34756 496 34812 524
rect 34876 496 34932 524
rect 34996 496 35052 524
rect 35116 496 35172 524
rect 35236 496 35292 524
rect 35356 496 35412 524
rect 35476 496 35532 524
rect 35596 496 35652 524
rect 35716 496 35772 524
rect 35836 496 35892 524
rect 35956 496 36012 524
rect 36076 496 36132 524
rect 36196 496 36252 524
rect 36316 496 36372 524
rect 36436 496 36492 524
rect 36556 496 36612 524
rect 36676 496 36732 524
rect 36796 496 36852 524
rect 36916 496 36972 524
rect 37036 496 37092 524
rect 37156 496 37212 524
rect 37276 496 37332 524
rect 37396 496 37452 524
rect 37516 496 37572 524
rect 37636 496 37692 524
rect 37756 496 37812 524
rect 37876 496 37932 524
rect 37996 496 38052 524
rect 38116 496 38172 524
rect 38236 496 38292 524
rect 38356 496 38412 524
rect 38476 496 38532 524
rect 38596 496 38652 524
rect 38716 496 38772 524
rect 38836 496 38892 524
rect 38956 496 39012 524
rect 39076 496 39132 524
rect 39196 496 39252 524
rect 39316 496 39372 524
rect 39436 496 39492 524
rect 39556 496 39612 524
rect 39676 496 39732 524
rect 39796 496 39852 524
rect 39916 496 39972 524
rect 40036 496 40092 524
rect 40156 496 40212 524
rect 40276 496 40332 524
rect 40396 496 40452 524
rect 40516 496 40572 524
rect 40636 496 40692 524
rect 40756 496 40812 524
rect 40876 496 40932 524
rect 40996 496 41052 524
rect 41116 496 41172 524
rect 41236 496 41292 524
rect 41356 496 41412 524
rect 41476 496 41532 524
rect 41596 496 41652 524
rect 41716 496 41772 524
rect 41836 496 41892 524
rect 41956 496 42012 524
rect 42076 496 42132 524
rect 42196 496 42252 524
rect 42316 496 42372 524
rect 42436 496 42492 524
rect 42556 496 42612 524
rect 42676 496 42732 524
rect 42796 496 42852 524
rect 42916 496 42972 524
rect 43036 496 43092 524
rect 43156 496 43212 524
rect 43276 496 43332 524
rect 43396 496 43452 524
rect 43516 496 43572 524
rect 43636 496 43692 524
rect 43756 496 43812 524
rect 43876 496 43932 524
rect 43996 496 44052 524
rect 44116 496 44172 524
rect 44236 496 44292 524
rect 44356 496 44412 524
rect 44476 496 44532 524
rect 44596 496 44652 524
rect 44716 496 44772 524
rect 44836 496 44892 524
rect 44956 496 45012 524
rect 45076 496 45132 524
rect 45196 496 45252 524
rect 45316 496 45372 524
rect 45436 496 45492 524
rect 45556 496 45612 524
rect 25848 -4328 25932 -4308
rect 25848 -4336 25868 -4328
rect 25876 -4336 25904 -4328
rect 25912 -4336 25932 -4328
rect 25968 -4328 26052 -4308
rect 25968 -4336 25988 -4328
rect 25996 -4336 26024 -4328
rect 26032 -4336 26052 -4328
rect 26088 -4328 26172 -4308
rect 26088 -4336 26108 -4328
rect 26116 -4336 26144 -4328
rect 26152 -4336 26172 -4328
rect 26208 -4328 26292 -4308
rect 26208 -4336 26228 -4328
rect 26236 -4336 26264 -4328
rect 26272 -4336 26292 -4328
rect 26328 -4328 26412 -4308
rect 26328 -4336 26348 -4328
rect 26356 -4336 26384 -4328
rect 26392 -4336 26412 -4328
rect 26448 -4328 26532 -4308
rect 26448 -4336 26468 -4328
rect 26476 -4336 26504 -4328
rect 26512 -4336 26532 -4328
rect 26568 -4328 26652 -4308
rect 26568 -4336 26588 -4328
rect 26596 -4336 26624 -4328
rect 26632 -4336 26652 -4328
rect 26688 -4328 26772 -4308
rect 26688 -4336 26708 -4328
rect 26716 -4336 26744 -4328
rect 26752 -4336 26772 -4328
rect 26808 -4328 26892 -4308
rect 26808 -4336 26828 -4328
rect 26836 -4336 26864 -4328
rect 26872 -4336 26892 -4328
rect 26928 -4328 27012 -4308
rect 26928 -4336 26948 -4328
rect 26956 -4336 26984 -4328
rect 26992 -4336 27012 -4328
rect 27048 -4328 27132 -4308
rect 27048 -4336 27068 -4328
rect 27076 -4336 27104 -4328
rect 27112 -4336 27132 -4328
rect 27168 -4328 27252 -4308
rect 27168 -4336 27188 -4328
rect 27196 -4336 27224 -4328
rect 27232 -4336 27252 -4328
rect 27288 -4328 27372 -4308
rect 27288 -4336 27308 -4328
rect 27316 -4336 27344 -4328
rect 27352 -4336 27372 -4328
rect 27408 -4328 27492 -4308
rect 27408 -4336 27428 -4328
rect 27436 -4336 27464 -4328
rect 27472 -4336 27492 -4328
rect 27528 -4328 27612 -4308
rect 27528 -4336 27548 -4328
rect 27556 -4336 27584 -4328
rect 27592 -4336 27612 -4328
rect 27648 -4328 27732 -4308
rect 27648 -4336 27668 -4328
rect 27676 -4336 27704 -4328
rect 27712 -4336 27732 -4328
rect 27768 -4328 27852 -4308
rect 27768 -4336 27788 -4328
rect 27796 -4336 27824 -4328
rect 27832 -4336 27852 -4328
rect 27888 -4328 27972 -4308
rect 27888 -4336 27908 -4328
rect 27916 -4336 27944 -4328
rect 27952 -4336 27972 -4328
rect 28008 -4328 28092 -4308
rect 28008 -4336 28028 -4328
rect 28036 -4336 28064 -4328
rect 28072 -4336 28092 -4328
rect 28128 -4328 28212 -4308
rect 28128 -4336 28148 -4328
rect 28156 -4336 28184 -4328
rect 28192 -4336 28212 -4328
rect 28248 -4328 28332 -4308
rect 28248 -4336 28268 -4328
rect 28276 -4336 28304 -4328
rect 28312 -4336 28332 -4328
rect 28368 -4328 28452 -4308
rect 28368 -4336 28388 -4328
rect 28396 -4336 28424 -4328
rect 28432 -4336 28452 -4328
rect 28488 -4328 28572 -4308
rect 28488 -4336 28508 -4328
rect 28516 -4336 28544 -4328
rect 28552 -4336 28572 -4328
rect 28608 -4328 28692 -4308
rect 28608 -4336 28628 -4328
rect 28636 -4336 28664 -4328
rect 28672 -4336 28692 -4328
rect 28728 -4328 28812 -4308
rect 28728 -4336 28748 -4328
rect 28756 -4336 28784 -4328
rect 28792 -4336 28812 -4328
rect 28848 -4328 28932 -4308
rect 28848 -4336 28868 -4328
rect 28876 -4336 28904 -4328
rect 28912 -4336 28932 -4328
rect 28968 -4328 29052 -4308
rect 28968 -4336 28988 -4328
rect 28996 -4336 29024 -4328
rect 29032 -4336 29052 -4328
rect 29088 -4328 29172 -4308
rect 29088 -4336 29108 -4328
rect 29116 -4336 29144 -4328
rect 29152 -4336 29172 -4328
rect 29208 -4328 29292 -4308
rect 29208 -4336 29228 -4328
rect 29236 -4336 29264 -4328
rect 29272 -4336 29292 -4328
rect 29328 -4328 29412 -4308
rect 29328 -4336 29348 -4328
rect 29356 -4336 29384 -4328
rect 29392 -4336 29412 -4328
rect 29448 -4328 29532 -4308
rect 29448 -4336 29468 -4328
rect 29476 -4336 29504 -4328
rect 29512 -4336 29532 -4328
rect 29568 -4328 29652 -4308
rect 29568 -4336 29588 -4328
rect 29596 -4336 29624 -4328
rect 29632 -4336 29652 -4328
rect 29688 -4328 29772 -4308
rect 29688 -4336 29708 -4328
rect 29716 -4336 29744 -4328
rect 29752 -4336 29772 -4328
rect 29808 -4328 29892 -4308
rect 29808 -4336 29828 -4328
rect 29836 -4336 29864 -4328
rect 29872 -4336 29892 -4328
rect 29928 -4328 30012 -4308
rect 29928 -4336 29948 -4328
rect 29956 -4336 29984 -4328
rect 29992 -4336 30012 -4328
rect 30048 -4328 30132 -4308
rect 30048 -4336 30068 -4328
rect 30076 -4336 30104 -4328
rect 30112 -4336 30132 -4328
rect 30168 -4328 30252 -4308
rect 30168 -4336 30188 -4328
rect 30196 -4336 30224 -4328
rect 30232 -4336 30252 -4328
rect 30288 -4328 30372 -4308
rect 30288 -4336 30308 -4328
rect 30316 -4336 30344 -4328
rect 30352 -4336 30372 -4328
rect 30408 -4328 30492 -4308
rect 30408 -4336 30428 -4328
rect 30436 -4336 30464 -4328
rect 30472 -4336 30492 -4328
rect 30528 -4328 30612 -4308
rect 30528 -4336 30548 -4328
rect 30556 -4336 30584 -4328
rect 30592 -4336 30612 -4328
rect 30648 -4328 30732 -4308
rect 30648 -4336 30668 -4328
rect 30676 -4336 30704 -4328
rect 30712 -4336 30732 -4328
rect 30768 -4328 30852 -4308
rect 30768 -4336 30788 -4328
rect 30796 -4336 30824 -4328
rect 30832 -4336 30852 -4328
rect 30888 -4328 30972 -4308
rect 30888 -4336 30908 -4328
rect 30916 -4336 30944 -4328
rect 30952 -4336 30972 -4328
rect 31008 -4328 31092 -4308
rect 31008 -4336 31028 -4328
rect 31036 -4336 31064 -4328
rect 31072 -4336 31092 -4328
rect 31128 -4328 31212 -4308
rect 31128 -4336 31148 -4328
rect 31156 -4336 31184 -4328
rect 31192 -4336 31212 -4328
rect 31248 -4328 31332 -4308
rect 31248 -4336 31268 -4328
rect 31276 -4336 31304 -4328
rect 31312 -4336 31332 -4328
rect 31368 -4328 31452 -4308
rect 31368 -4336 31388 -4328
rect 31396 -4336 31424 -4328
rect 31432 -4336 31452 -4328
rect 31488 -4328 31572 -4308
rect 31488 -4336 31508 -4328
rect 31516 -4336 31544 -4328
rect 31552 -4336 31572 -4328
rect 31608 -4328 31692 -4308
rect 31608 -4336 31628 -4328
rect 31636 -4336 31664 -4328
rect 31672 -4336 31692 -4328
rect 31728 -4328 31812 -4308
rect 31728 -4336 31748 -4328
rect 31756 -4336 31784 -4328
rect 31792 -4336 31812 -4328
rect 31848 -4328 31932 -4308
rect 31848 -4336 31868 -4328
rect 31876 -4336 31904 -4328
rect 31912 -4336 31932 -4328
rect 31968 -4328 32052 -4308
rect 31968 -4336 31988 -4328
rect 31996 -4336 32024 -4328
rect 32032 -4336 32052 -4328
rect 32088 -4328 32172 -4308
rect 32088 -4336 32108 -4328
rect 32116 -4336 32144 -4328
rect 32152 -4336 32172 -4328
rect 32208 -4328 32292 -4308
rect 32208 -4336 32228 -4328
rect 32236 -4336 32264 -4328
rect 32272 -4336 32292 -4328
rect 32328 -4328 32412 -4308
rect 32328 -4336 32348 -4328
rect 32356 -4336 32384 -4328
rect 32392 -4336 32412 -4328
rect 32448 -4328 32532 -4308
rect 32448 -4336 32468 -4328
rect 32476 -4336 32504 -4328
rect 32512 -4336 32532 -4328
rect 32568 -4328 32652 -4308
rect 32568 -4336 32588 -4328
rect 32596 -4336 32624 -4328
rect 32632 -4336 32652 -4328
rect 32688 -4328 32772 -4308
rect 32688 -4336 32708 -4328
rect 32716 -4336 32744 -4328
rect 32752 -4336 32772 -4328
rect 32808 -4328 32892 -4308
rect 32808 -4336 32828 -4328
rect 32836 -4336 32864 -4328
rect 32872 -4336 32892 -4328
rect 32928 -4328 33012 -4308
rect 32928 -4336 32948 -4328
rect 32956 -4336 32984 -4328
rect 32992 -4336 33012 -4328
rect 33048 -4328 33132 -4308
rect 33048 -4336 33068 -4328
rect 33076 -4336 33104 -4328
rect 33112 -4336 33132 -4328
rect 33168 -4328 33252 -4308
rect 33168 -4336 33188 -4328
rect 33196 -4336 33224 -4328
rect 33232 -4336 33252 -4328
rect 33288 -4328 33372 -4308
rect 33288 -4336 33308 -4328
rect 33316 -4336 33344 -4328
rect 33352 -4336 33372 -4328
rect 33408 -4328 33492 -4308
rect 33408 -4336 33428 -4328
rect 33436 -4336 33464 -4328
rect 33472 -4336 33492 -4328
rect 33528 -4328 33612 -4308
rect 33528 -4336 33548 -4328
rect 33556 -4336 33584 -4328
rect 33592 -4336 33612 -4328
rect 33648 -4328 33732 -4308
rect 33648 -4336 33668 -4328
rect 33676 -4336 33704 -4328
rect 33712 -4336 33732 -4328
rect 33768 -4328 33852 -4308
rect 33768 -4336 33788 -4328
rect 33796 -4336 33824 -4328
rect 33832 -4336 33852 -4328
rect 33888 -4328 33972 -4308
rect 33888 -4336 33908 -4328
rect 33916 -4336 33944 -4328
rect 33952 -4336 33972 -4328
rect 34008 -4328 34092 -4308
rect 34008 -4336 34028 -4328
rect 34036 -4336 34064 -4328
rect 34072 -4336 34092 -4328
rect 34128 -4328 34212 -4308
rect 34128 -4336 34148 -4328
rect 34156 -4336 34184 -4328
rect 34192 -4336 34212 -4328
rect 34248 -4328 34332 -4308
rect 34248 -4336 34268 -4328
rect 34276 -4336 34304 -4328
rect 34312 -4336 34332 -4328
rect 34368 -4328 34452 -4308
rect 34368 -4336 34388 -4328
rect 34396 -4336 34424 -4328
rect 34432 -4336 34452 -4328
rect 34488 -4328 34572 -4308
rect 34488 -4336 34508 -4328
rect 34516 -4336 34544 -4328
rect 34552 -4336 34572 -4328
rect 34608 -4328 34692 -4308
rect 34608 -4336 34628 -4328
rect 34636 -4336 34664 -4328
rect 34672 -4336 34692 -4328
rect 34728 -4328 34812 -4308
rect 34728 -4336 34748 -4328
rect 34756 -4336 34784 -4328
rect 34792 -4336 34812 -4328
rect 34848 -4328 34932 -4308
rect 34848 -4336 34868 -4328
rect 34876 -4336 34904 -4328
rect 34912 -4336 34932 -4328
rect 34968 -4328 35052 -4308
rect 34968 -4336 34988 -4328
rect 34996 -4336 35024 -4328
rect 35032 -4336 35052 -4328
rect 35088 -4328 35172 -4308
rect 35088 -4336 35108 -4328
rect 35116 -4336 35144 -4328
rect 35152 -4336 35172 -4328
rect 35208 -4328 35292 -4308
rect 35208 -4336 35228 -4328
rect 35236 -4336 35264 -4328
rect 35272 -4336 35292 -4328
rect 35328 -4328 35412 -4308
rect 35328 -4336 35348 -4328
rect 35356 -4336 35384 -4328
rect 35392 -4336 35412 -4328
rect 35448 -4328 35532 -4308
rect 35448 -4336 35468 -4328
rect 35476 -4336 35504 -4328
rect 35512 -4336 35532 -4328
rect 35568 -4328 35652 -4308
rect 35568 -4336 35588 -4328
rect 35596 -4336 35624 -4328
rect 35632 -4336 35652 -4328
rect 35688 -4328 35772 -4308
rect 35688 -4336 35708 -4328
rect 35716 -4336 35744 -4328
rect 35752 -4336 35772 -4328
rect 35808 -4328 35892 -4308
rect 35808 -4336 35828 -4328
rect 35836 -4336 35864 -4328
rect 35872 -4336 35892 -4328
rect 35928 -4328 36012 -4308
rect 35928 -4336 35948 -4328
rect 35956 -4336 35984 -4328
rect 35992 -4336 36012 -4328
rect 36048 -4328 36132 -4308
rect 36048 -4336 36068 -4328
rect 36076 -4336 36104 -4328
rect 36112 -4336 36132 -4328
rect 36168 -4328 36252 -4308
rect 36168 -4336 36188 -4328
rect 36196 -4336 36224 -4328
rect 36232 -4336 36252 -4328
rect 36288 -4328 36372 -4308
rect 36288 -4336 36308 -4328
rect 36316 -4336 36344 -4328
rect 36352 -4336 36372 -4328
rect 36408 -4328 36492 -4308
rect 36408 -4336 36428 -4328
rect 36436 -4336 36464 -4328
rect 36472 -4336 36492 -4328
rect 36528 -4328 36612 -4308
rect 36528 -4336 36548 -4328
rect 36556 -4336 36584 -4328
rect 36592 -4336 36612 -4328
rect 36648 -4328 36732 -4308
rect 36648 -4336 36668 -4328
rect 36676 -4336 36704 -4328
rect 36712 -4336 36732 -4328
rect 36768 -4328 36852 -4308
rect 36768 -4336 36788 -4328
rect 36796 -4336 36824 -4328
rect 36832 -4336 36852 -4328
rect 36888 -4328 36972 -4308
rect 36888 -4336 36908 -4328
rect 36916 -4336 36944 -4328
rect 36952 -4336 36972 -4328
rect 37008 -4328 37092 -4308
rect 37008 -4336 37028 -4328
rect 37036 -4336 37064 -4328
rect 37072 -4336 37092 -4328
rect 37128 -4328 37212 -4308
rect 37128 -4336 37148 -4328
rect 37156 -4336 37184 -4328
rect 37192 -4336 37212 -4328
rect 37248 -4328 37332 -4308
rect 37248 -4336 37268 -4328
rect 37276 -4336 37304 -4328
rect 37312 -4336 37332 -4328
rect 37368 -4328 37452 -4308
rect 37368 -4336 37388 -4328
rect 37396 -4336 37424 -4328
rect 37432 -4336 37452 -4328
rect 37488 -4328 37572 -4308
rect 37488 -4336 37508 -4328
rect 37516 -4336 37544 -4328
rect 37552 -4336 37572 -4328
rect 37608 -4328 37692 -4308
rect 37608 -4336 37628 -4328
rect 37636 -4336 37664 -4328
rect 37672 -4336 37692 -4328
rect 37728 -4328 37812 -4308
rect 37728 -4336 37748 -4328
rect 37756 -4336 37784 -4328
rect 37792 -4336 37812 -4328
rect 37848 -4328 37932 -4308
rect 37848 -4336 37868 -4328
rect 37876 -4336 37904 -4328
rect 37912 -4336 37932 -4328
rect 37968 -4328 38052 -4308
rect 37968 -4336 37988 -4328
rect 37996 -4336 38024 -4328
rect 38032 -4336 38052 -4328
rect 38088 -4328 38172 -4308
rect 38088 -4336 38108 -4328
rect 38116 -4336 38144 -4328
rect 38152 -4336 38172 -4328
rect 38208 -4328 38292 -4308
rect 38208 -4336 38228 -4328
rect 38236 -4336 38264 -4328
rect 38272 -4336 38292 -4328
rect 38328 -4328 38412 -4308
rect 38328 -4336 38348 -4328
rect 38356 -4336 38384 -4328
rect 38392 -4336 38412 -4328
rect 38448 -4328 38532 -4308
rect 38448 -4336 38468 -4328
rect 38476 -4336 38504 -4328
rect 38512 -4336 38532 -4328
rect 38568 -4328 38652 -4308
rect 38568 -4336 38588 -4328
rect 38596 -4336 38624 -4328
rect 38632 -4336 38652 -4328
rect 38688 -4328 38772 -4308
rect 38688 -4336 38708 -4328
rect 38716 -4336 38744 -4328
rect 38752 -4336 38772 -4328
rect 38808 -4328 38892 -4308
rect 38808 -4336 38828 -4328
rect 38836 -4336 38864 -4328
rect 38872 -4336 38892 -4328
rect 38928 -4328 39012 -4308
rect 38928 -4336 38948 -4328
rect 38956 -4336 38984 -4328
rect 38992 -4336 39012 -4328
rect 39048 -4328 39132 -4308
rect 39048 -4336 39068 -4328
rect 39076 -4336 39104 -4328
rect 39112 -4336 39132 -4328
rect 39168 -4328 39252 -4308
rect 39168 -4336 39188 -4328
rect 39196 -4336 39224 -4328
rect 39232 -4336 39252 -4328
rect 39288 -4328 39372 -4308
rect 39288 -4336 39308 -4328
rect 39316 -4336 39344 -4328
rect 39352 -4336 39372 -4328
rect 39408 -4328 39492 -4308
rect 39408 -4336 39428 -4328
rect 39436 -4336 39464 -4328
rect 39472 -4336 39492 -4328
rect 39528 -4328 39612 -4308
rect 39528 -4336 39548 -4328
rect 39556 -4336 39584 -4328
rect 39592 -4336 39612 -4328
rect 39648 -4328 39732 -4308
rect 39648 -4336 39668 -4328
rect 39676 -4336 39704 -4328
rect 39712 -4336 39732 -4328
rect 39768 -4328 39852 -4308
rect 39768 -4336 39788 -4328
rect 39796 -4336 39824 -4328
rect 39832 -4336 39852 -4328
rect 39888 -4328 39972 -4308
rect 39888 -4336 39908 -4328
rect 39916 -4336 39944 -4328
rect 39952 -4336 39972 -4328
rect 40008 -4328 40092 -4308
rect 40008 -4336 40028 -4328
rect 40036 -4336 40064 -4328
rect 40072 -4336 40092 -4328
rect 40128 -4328 40212 -4308
rect 40128 -4336 40148 -4328
rect 40156 -4336 40184 -4328
rect 40192 -4336 40212 -4328
rect 40248 -4328 40332 -4308
rect 40248 -4336 40268 -4328
rect 40276 -4336 40304 -4328
rect 40312 -4336 40332 -4328
rect 40368 -4328 40452 -4308
rect 40368 -4336 40388 -4328
rect 40396 -4336 40424 -4328
rect 40432 -4336 40452 -4328
rect 40488 -4328 40572 -4308
rect 40488 -4336 40508 -4328
rect 40516 -4336 40544 -4328
rect 40552 -4336 40572 -4328
rect 40608 -4328 40692 -4308
rect 40608 -4336 40628 -4328
rect 40636 -4336 40664 -4328
rect 40672 -4336 40692 -4328
rect 40728 -4328 40812 -4308
rect 40728 -4336 40748 -4328
rect 40756 -4336 40784 -4328
rect 40792 -4336 40812 -4328
rect 40848 -4328 40932 -4308
rect 40848 -4336 40868 -4328
rect 40876 -4336 40904 -4328
rect 40912 -4336 40932 -4328
rect 40968 -4328 41052 -4308
rect 40968 -4336 40988 -4328
rect 40996 -4336 41024 -4328
rect 41032 -4336 41052 -4328
rect 41088 -4328 41172 -4308
rect 41088 -4336 41108 -4328
rect 41116 -4336 41144 -4328
rect 41152 -4336 41172 -4328
rect 41208 -4328 41292 -4308
rect 41208 -4336 41228 -4328
rect 41236 -4336 41264 -4328
rect 41272 -4336 41292 -4328
rect 41328 -4328 41412 -4308
rect 41328 -4336 41348 -4328
rect 41356 -4336 41384 -4328
rect 41392 -4336 41412 -4328
rect 41448 -4328 41532 -4308
rect 41448 -4336 41468 -4328
rect 41476 -4336 41504 -4328
rect 41512 -4336 41532 -4328
rect 41568 -4328 41652 -4308
rect 41568 -4336 41588 -4328
rect 41596 -4336 41624 -4328
rect 41632 -4336 41652 -4328
rect 41688 -4328 41772 -4308
rect 41688 -4336 41708 -4328
rect 41716 -4336 41744 -4328
rect 41752 -4336 41772 -4328
rect 41808 -4328 41892 -4308
rect 41808 -4336 41828 -4328
rect 41836 -4336 41864 -4328
rect 41872 -4336 41892 -4328
rect 41928 -4328 42012 -4308
rect 41928 -4336 41948 -4328
rect 41956 -4336 41984 -4328
rect 41992 -4336 42012 -4328
rect 42048 -4328 42132 -4308
rect 42048 -4336 42068 -4328
rect 42076 -4336 42104 -4328
rect 42112 -4336 42132 -4328
rect 42168 -4328 42252 -4308
rect 42168 -4336 42188 -4328
rect 42196 -4336 42224 -4328
rect 42232 -4336 42252 -4328
rect 42288 -4328 42372 -4308
rect 42288 -4336 42308 -4328
rect 42316 -4336 42344 -4328
rect 42352 -4336 42372 -4328
rect 42408 -4328 42492 -4308
rect 42408 -4336 42428 -4328
rect 42436 -4336 42464 -4328
rect 42472 -4336 42492 -4328
rect 42528 -4328 42612 -4308
rect 42528 -4336 42548 -4328
rect 42556 -4336 42584 -4328
rect 42592 -4336 42612 -4328
rect 42648 -4328 42732 -4308
rect 42648 -4336 42668 -4328
rect 42676 -4336 42704 -4328
rect 42712 -4336 42732 -4328
rect 42768 -4328 42852 -4308
rect 42768 -4336 42788 -4328
rect 42796 -4336 42824 -4328
rect 42832 -4336 42852 -4328
rect 42888 -4328 42972 -4308
rect 42888 -4336 42908 -4328
rect 42916 -4336 42944 -4328
rect 42952 -4336 42972 -4328
rect 43008 -4328 43092 -4308
rect 43008 -4336 43028 -4328
rect 43036 -4336 43064 -4328
rect 43072 -4336 43092 -4328
rect 43128 -4328 43212 -4308
rect 43128 -4336 43148 -4328
rect 43156 -4336 43184 -4328
rect 43192 -4336 43212 -4328
rect 43248 -4328 43332 -4308
rect 43248 -4336 43268 -4328
rect 43276 -4336 43304 -4328
rect 43312 -4336 43332 -4328
rect 43368 -4328 43452 -4308
rect 43368 -4336 43388 -4328
rect 43396 -4336 43424 -4328
rect 43432 -4336 43452 -4328
rect 43488 -4328 43572 -4308
rect 43488 -4336 43508 -4328
rect 43516 -4336 43544 -4328
rect 43552 -4336 43572 -4328
rect 43608 -4328 43692 -4308
rect 43608 -4336 43628 -4328
rect 43636 -4336 43664 -4328
rect 43672 -4336 43692 -4328
rect 43728 -4328 43812 -4308
rect 43728 -4336 43748 -4328
rect 43756 -4336 43784 -4328
rect 43792 -4336 43812 -4328
rect 43848 -4328 43932 -4308
rect 43848 -4336 43868 -4328
rect 43876 -4336 43904 -4328
rect 43912 -4336 43932 -4328
rect 43968 -4328 44052 -4308
rect 43968 -4336 43988 -4328
rect 43996 -4336 44024 -4328
rect 44032 -4336 44052 -4328
rect 44088 -4328 44172 -4308
rect 44088 -4336 44108 -4328
rect 44116 -4336 44144 -4328
rect 44152 -4336 44172 -4328
rect 44208 -4328 44292 -4308
rect 44208 -4336 44228 -4328
rect 44236 -4336 44264 -4328
rect 44272 -4336 44292 -4328
rect 44328 -4328 44412 -4308
rect 44328 -4336 44348 -4328
rect 44356 -4336 44384 -4328
rect 44392 -4336 44412 -4328
rect 44448 -4328 44532 -4308
rect 44448 -4336 44468 -4328
rect 44476 -4336 44504 -4328
rect 44512 -4336 44532 -4328
rect 44568 -4328 44652 -4308
rect 44568 -4336 44588 -4328
rect 44596 -4336 44624 -4328
rect 44632 -4336 44652 -4328
rect 44688 -4328 44772 -4308
rect 44688 -4336 44708 -4328
rect 44716 -4336 44744 -4328
rect 44752 -4336 44772 -4328
rect 44808 -4328 44892 -4308
rect 44808 -4336 44828 -4328
rect 44836 -4336 44864 -4328
rect 44872 -4336 44892 -4328
rect 44928 -4328 45012 -4308
rect 44928 -4336 44948 -4328
rect 44956 -4336 44984 -4328
rect 44992 -4336 45012 -4328
rect 45048 -4328 45132 -4308
rect 45048 -4336 45068 -4328
rect 45076 -4336 45104 -4328
rect 45112 -4336 45132 -4328
rect 45168 -4328 45252 -4308
rect 45168 -4336 45188 -4328
rect 45196 -4336 45224 -4328
rect 45232 -4336 45252 -4328
rect 45288 -4328 45372 -4308
rect 45288 -4336 45308 -4328
rect 45316 -4336 45344 -4328
rect 45352 -4336 45372 -4328
rect 45408 -4328 45492 -4308
rect 45408 -4336 45428 -4328
rect 45436 -4336 45464 -4328
rect 45472 -4336 45492 -4328
rect 45528 -4328 45612 -4308
rect 45528 -4336 45548 -4328
rect 45556 -4336 45584 -4328
rect 45592 -4336 45612 -4328
rect 25876 -4364 25932 -4336
rect 25996 -4364 26052 -4336
rect 26116 -4364 26172 -4336
rect 26236 -4364 26292 -4336
rect 26356 -4364 26412 -4336
rect 26476 -4364 26532 -4336
rect 26596 -4364 26652 -4336
rect 26716 -4364 26772 -4336
rect 26836 -4364 26892 -4336
rect 26956 -4364 27012 -4336
rect 27076 -4364 27132 -4336
rect 27196 -4364 27252 -4336
rect 27316 -4364 27372 -4336
rect 27436 -4364 27492 -4336
rect 27556 -4364 27612 -4336
rect 27676 -4364 27732 -4336
rect 27796 -4364 27852 -4336
rect 27916 -4364 27972 -4336
rect 28036 -4364 28092 -4336
rect 28156 -4364 28212 -4336
rect 28276 -4364 28332 -4336
rect 28396 -4364 28452 -4336
rect 28516 -4364 28572 -4336
rect 28636 -4364 28692 -4336
rect 28756 -4364 28812 -4336
rect 28876 -4364 28932 -4336
rect 28996 -4364 29052 -4336
rect 29116 -4364 29172 -4336
rect 29236 -4364 29292 -4336
rect 29356 -4364 29412 -4336
rect 29476 -4364 29532 -4336
rect 29596 -4364 29652 -4336
rect 29716 -4364 29772 -4336
rect 29836 -4364 29892 -4336
rect 29956 -4364 30012 -4336
rect 30076 -4364 30132 -4336
rect 30196 -4364 30252 -4336
rect 30316 -4364 30372 -4336
rect 30436 -4364 30492 -4336
rect 30556 -4364 30612 -4336
rect 30676 -4364 30732 -4336
rect 30796 -4364 30852 -4336
rect 30916 -4364 30972 -4336
rect 31036 -4364 31092 -4336
rect 31156 -4364 31212 -4336
rect 31276 -4364 31332 -4336
rect 31396 -4364 31452 -4336
rect 31516 -4364 31572 -4336
rect 31636 -4364 31692 -4336
rect 31756 -4364 31812 -4336
rect 31876 -4364 31932 -4336
rect 31996 -4364 32052 -4336
rect 32116 -4364 32172 -4336
rect 32236 -4364 32292 -4336
rect 32356 -4364 32412 -4336
rect 32476 -4364 32532 -4336
rect 32596 -4364 32652 -4336
rect 32716 -4364 32772 -4336
rect 32836 -4364 32892 -4336
rect 32956 -4364 33012 -4336
rect 33076 -4364 33132 -4336
rect 33196 -4364 33252 -4336
rect 33316 -4364 33372 -4336
rect 33436 -4364 33492 -4336
rect 33556 -4364 33612 -4336
rect 33676 -4364 33732 -4336
rect 33796 -4364 33852 -4336
rect 33916 -4364 33972 -4336
rect 34036 -4364 34092 -4336
rect 34156 -4364 34212 -4336
rect 34276 -4364 34332 -4336
rect 34396 -4364 34452 -4336
rect 34516 -4364 34572 -4336
rect 34636 -4364 34692 -4336
rect 34756 -4364 34812 -4336
rect 34876 -4364 34932 -4336
rect 34996 -4364 35052 -4336
rect 35116 -4364 35172 -4336
rect 35236 -4364 35292 -4336
rect 35356 -4364 35412 -4336
rect 35476 -4364 35532 -4336
rect 35596 -4364 35652 -4336
rect 35716 -4364 35772 -4336
rect 35836 -4364 35892 -4336
rect 35956 -4364 36012 -4336
rect 36076 -4364 36132 -4336
rect 36196 -4364 36252 -4336
rect 36316 -4364 36372 -4336
rect 36436 -4364 36492 -4336
rect 36556 -4364 36612 -4336
rect 36676 -4364 36732 -4336
rect 36796 -4364 36852 -4336
rect 36916 -4364 36972 -4336
rect 37036 -4364 37092 -4336
rect 37156 -4364 37212 -4336
rect 37276 -4364 37332 -4336
rect 37396 -4364 37452 -4336
rect 37516 -4364 37572 -4336
rect 37636 -4364 37692 -4336
rect 37756 -4364 37812 -4336
rect 37876 -4364 37932 -4336
rect 37996 -4364 38052 -4336
rect 38116 -4364 38172 -4336
rect 38236 -4364 38292 -4336
rect 38356 -4364 38412 -4336
rect 38476 -4364 38532 -4336
rect 38596 -4364 38652 -4336
rect 38716 -4364 38772 -4336
rect 38836 -4364 38892 -4336
rect 38956 -4364 39012 -4336
rect 39076 -4364 39132 -4336
rect 39196 -4364 39252 -4336
rect 39316 -4364 39372 -4336
rect 39436 -4364 39492 -4336
rect 39556 -4364 39612 -4336
rect 39676 -4364 39732 -4336
rect 39796 -4364 39852 -4336
rect 39916 -4364 39972 -4336
rect 40036 -4364 40092 -4336
rect 40156 -4364 40212 -4336
rect 40276 -4364 40332 -4336
rect 40396 -4364 40452 -4336
rect 40516 -4364 40572 -4336
rect 40636 -4364 40692 -4336
rect 40756 -4364 40812 -4336
rect 40876 -4364 40932 -4336
rect 40996 -4364 41052 -4336
rect 41116 -4364 41172 -4336
rect 41236 -4364 41292 -4336
rect 41356 -4364 41412 -4336
rect 41476 -4364 41532 -4336
rect 41596 -4364 41652 -4336
rect 41716 -4364 41772 -4336
rect 41836 -4364 41892 -4336
rect 41956 -4364 42012 -4336
rect 42076 -4364 42132 -4336
rect 42196 -4364 42252 -4336
rect 42316 -4364 42372 -4336
rect 42436 -4364 42492 -4336
rect 42556 -4364 42612 -4336
rect 42676 -4364 42732 -4336
rect 42796 -4364 42852 -4336
rect 42916 -4364 42972 -4336
rect 43036 -4364 43092 -4336
rect 43156 -4364 43212 -4336
rect 43276 -4364 43332 -4336
rect 43396 -4364 43452 -4336
rect 43516 -4364 43572 -4336
rect 43636 -4364 43692 -4336
rect 43756 -4364 43812 -4336
rect 43876 -4364 43932 -4336
rect 43996 -4364 44052 -4336
rect 44116 -4364 44172 -4336
rect 44236 -4364 44292 -4336
rect 44356 -4364 44412 -4336
rect 44476 -4364 44532 -4336
rect 44596 -4364 44652 -4336
rect 44716 -4364 44772 -4336
rect 44836 -4364 44892 -4336
rect 44956 -4364 45012 -4336
rect 45076 -4364 45132 -4336
rect 45196 -4364 45252 -4336
rect 45316 -4364 45372 -4336
rect 45436 -4364 45492 -4336
rect 45556 -4364 45612 -4336
rect 25848 -4508 25932 -4488
rect 25848 -4516 25868 -4508
rect 25876 -4516 25904 -4508
rect 25912 -4516 25932 -4508
rect 25968 -4508 26052 -4488
rect 25968 -4516 25988 -4508
rect 25996 -4516 26024 -4508
rect 26032 -4516 26052 -4508
rect 26088 -4508 26172 -4488
rect 26088 -4516 26108 -4508
rect 26116 -4516 26144 -4508
rect 26152 -4516 26172 -4508
rect 26208 -4508 26292 -4488
rect 26208 -4516 26228 -4508
rect 26236 -4516 26264 -4508
rect 26272 -4516 26292 -4508
rect 26328 -4508 26412 -4488
rect 26328 -4516 26348 -4508
rect 26356 -4516 26384 -4508
rect 26392 -4516 26412 -4508
rect 26448 -4508 26532 -4488
rect 26448 -4516 26468 -4508
rect 26476 -4516 26504 -4508
rect 26512 -4516 26532 -4508
rect 26568 -4508 26652 -4488
rect 26568 -4516 26588 -4508
rect 26596 -4516 26624 -4508
rect 26632 -4516 26652 -4508
rect 26688 -4508 26772 -4488
rect 26688 -4516 26708 -4508
rect 26716 -4516 26744 -4508
rect 26752 -4516 26772 -4508
rect 26808 -4508 26892 -4488
rect 26808 -4516 26828 -4508
rect 26836 -4516 26864 -4508
rect 26872 -4516 26892 -4508
rect 26928 -4508 27012 -4488
rect 26928 -4516 26948 -4508
rect 26956 -4516 26984 -4508
rect 26992 -4516 27012 -4508
rect 27048 -4508 27132 -4488
rect 27048 -4516 27068 -4508
rect 27076 -4516 27104 -4508
rect 27112 -4516 27132 -4508
rect 27168 -4508 27252 -4488
rect 27168 -4516 27188 -4508
rect 27196 -4516 27224 -4508
rect 27232 -4516 27252 -4508
rect 27288 -4508 27372 -4488
rect 27288 -4516 27308 -4508
rect 27316 -4516 27344 -4508
rect 27352 -4516 27372 -4508
rect 27408 -4508 27492 -4488
rect 27408 -4516 27428 -4508
rect 27436 -4516 27464 -4508
rect 27472 -4516 27492 -4508
rect 27528 -4508 27612 -4488
rect 27528 -4516 27548 -4508
rect 27556 -4516 27584 -4508
rect 27592 -4516 27612 -4508
rect 27648 -4508 27732 -4488
rect 27648 -4516 27668 -4508
rect 27676 -4516 27704 -4508
rect 27712 -4516 27732 -4508
rect 27768 -4508 27852 -4488
rect 27768 -4516 27788 -4508
rect 27796 -4516 27824 -4508
rect 27832 -4516 27852 -4508
rect 27888 -4508 27972 -4488
rect 27888 -4516 27908 -4508
rect 27916 -4516 27944 -4508
rect 27952 -4516 27972 -4508
rect 28008 -4508 28092 -4488
rect 28008 -4516 28028 -4508
rect 28036 -4516 28064 -4508
rect 28072 -4516 28092 -4508
rect 28128 -4508 28212 -4488
rect 28128 -4516 28148 -4508
rect 28156 -4516 28184 -4508
rect 28192 -4516 28212 -4508
rect 28248 -4508 28332 -4488
rect 28248 -4516 28268 -4508
rect 28276 -4516 28304 -4508
rect 28312 -4516 28332 -4508
rect 28368 -4508 28452 -4488
rect 28368 -4516 28388 -4508
rect 28396 -4516 28424 -4508
rect 28432 -4516 28452 -4508
rect 28488 -4508 28572 -4488
rect 28488 -4516 28508 -4508
rect 28516 -4516 28544 -4508
rect 28552 -4516 28572 -4508
rect 28608 -4508 28692 -4488
rect 28608 -4516 28628 -4508
rect 28636 -4516 28664 -4508
rect 28672 -4516 28692 -4508
rect 28728 -4508 28812 -4488
rect 28728 -4516 28748 -4508
rect 28756 -4516 28784 -4508
rect 28792 -4516 28812 -4508
rect 28848 -4508 28932 -4488
rect 28848 -4516 28868 -4508
rect 28876 -4516 28904 -4508
rect 28912 -4516 28932 -4508
rect 28968 -4508 29052 -4488
rect 28968 -4516 28988 -4508
rect 28996 -4516 29024 -4508
rect 29032 -4516 29052 -4508
rect 29088 -4508 29172 -4488
rect 29088 -4516 29108 -4508
rect 29116 -4516 29144 -4508
rect 29152 -4516 29172 -4508
rect 29208 -4508 29292 -4488
rect 29208 -4516 29228 -4508
rect 29236 -4516 29264 -4508
rect 29272 -4516 29292 -4508
rect 29328 -4508 29412 -4488
rect 29328 -4516 29348 -4508
rect 29356 -4516 29384 -4508
rect 29392 -4516 29412 -4508
rect 29448 -4508 29532 -4488
rect 29448 -4516 29468 -4508
rect 29476 -4516 29504 -4508
rect 29512 -4516 29532 -4508
rect 29568 -4508 29652 -4488
rect 29568 -4516 29588 -4508
rect 29596 -4516 29624 -4508
rect 29632 -4516 29652 -4508
rect 29688 -4508 29772 -4488
rect 29688 -4516 29708 -4508
rect 29716 -4516 29744 -4508
rect 29752 -4516 29772 -4508
rect 29808 -4508 29892 -4488
rect 29808 -4516 29828 -4508
rect 29836 -4516 29864 -4508
rect 29872 -4516 29892 -4508
rect 29928 -4508 30012 -4488
rect 29928 -4516 29948 -4508
rect 29956 -4516 29984 -4508
rect 29992 -4516 30012 -4508
rect 30048 -4508 30132 -4488
rect 30048 -4516 30068 -4508
rect 30076 -4516 30104 -4508
rect 30112 -4516 30132 -4508
rect 30168 -4508 30252 -4488
rect 30168 -4516 30188 -4508
rect 30196 -4516 30224 -4508
rect 30232 -4516 30252 -4508
rect 30288 -4508 30372 -4488
rect 30288 -4516 30308 -4508
rect 30316 -4516 30344 -4508
rect 30352 -4516 30372 -4508
rect 30408 -4508 30492 -4488
rect 30408 -4516 30428 -4508
rect 30436 -4516 30464 -4508
rect 30472 -4516 30492 -4508
rect 30528 -4508 30612 -4488
rect 30528 -4516 30548 -4508
rect 30556 -4516 30584 -4508
rect 30592 -4516 30612 -4508
rect 30648 -4508 30732 -4488
rect 30648 -4516 30668 -4508
rect 30676 -4516 30704 -4508
rect 30712 -4516 30732 -4508
rect 30768 -4508 30852 -4488
rect 30768 -4516 30788 -4508
rect 30796 -4516 30824 -4508
rect 30832 -4516 30852 -4508
rect 30888 -4508 30972 -4488
rect 30888 -4516 30908 -4508
rect 30916 -4516 30944 -4508
rect 30952 -4516 30972 -4508
rect 31008 -4508 31092 -4488
rect 31008 -4516 31028 -4508
rect 31036 -4516 31064 -4508
rect 31072 -4516 31092 -4508
rect 31128 -4508 31212 -4488
rect 31128 -4516 31148 -4508
rect 31156 -4516 31184 -4508
rect 31192 -4516 31212 -4508
rect 31248 -4508 31332 -4488
rect 31248 -4516 31268 -4508
rect 31276 -4516 31304 -4508
rect 31312 -4516 31332 -4508
rect 31368 -4508 31452 -4488
rect 31368 -4516 31388 -4508
rect 31396 -4516 31424 -4508
rect 31432 -4516 31452 -4508
rect 31488 -4508 31572 -4488
rect 31488 -4516 31508 -4508
rect 31516 -4516 31544 -4508
rect 31552 -4516 31572 -4508
rect 31608 -4508 31692 -4488
rect 31608 -4516 31628 -4508
rect 31636 -4516 31664 -4508
rect 31672 -4516 31692 -4508
rect 31728 -4508 31812 -4488
rect 31728 -4516 31748 -4508
rect 31756 -4516 31784 -4508
rect 31792 -4516 31812 -4508
rect 31848 -4508 31932 -4488
rect 31848 -4516 31868 -4508
rect 31876 -4516 31904 -4508
rect 31912 -4516 31932 -4508
rect 31968 -4508 32052 -4488
rect 31968 -4516 31988 -4508
rect 31996 -4516 32024 -4508
rect 32032 -4516 32052 -4508
rect 32088 -4508 32172 -4488
rect 32088 -4516 32108 -4508
rect 32116 -4516 32144 -4508
rect 32152 -4516 32172 -4508
rect 32208 -4508 32292 -4488
rect 32208 -4516 32228 -4508
rect 32236 -4516 32264 -4508
rect 32272 -4516 32292 -4508
rect 32328 -4508 32412 -4488
rect 32328 -4516 32348 -4508
rect 32356 -4516 32384 -4508
rect 32392 -4516 32412 -4508
rect 32448 -4508 32532 -4488
rect 32448 -4516 32468 -4508
rect 32476 -4516 32504 -4508
rect 32512 -4516 32532 -4508
rect 32568 -4508 32652 -4488
rect 32568 -4516 32588 -4508
rect 32596 -4516 32624 -4508
rect 32632 -4516 32652 -4508
rect 32688 -4508 32772 -4488
rect 32688 -4516 32708 -4508
rect 32716 -4516 32744 -4508
rect 32752 -4516 32772 -4508
rect 32808 -4508 32892 -4488
rect 32808 -4516 32828 -4508
rect 32836 -4516 32864 -4508
rect 32872 -4516 32892 -4508
rect 32928 -4508 33012 -4488
rect 32928 -4516 32948 -4508
rect 32956 -4516 32984 -4508
rect 32992 -4516 33012 -4508
rect 33048 -4508 33132 -4488
rect 33048 -4516 33068 -4508
rect 33076 -4516 33104 -4508
rect 33112 -4516 33132 -4508
rect 33168 -4508 33252 -4488
rect 33168 -4516 33188 -4508
rect 33196 -4516 33224 -4508
rect 33232 -4516 33252 -4508
rect 33288 -4508 33372 -4488
rect 33288 -4516 33308 -4508
rect 33316 -4516 33344 -4508
rect 33352 -4516 33372 -4508
rect 33408 -4508 33492 -4488
rect 33408 -4516 33428 -4508
rect 33436 -4516 33464 -4508
rect 33472 -4516 33492 -4508
rect 33528 -4508 33612 -4488
rect 33528 -4516 33548 -4508
rect 33556 -4516 33584 -4508
rect 33592 -4516 33612 -4508
rect 33648 -4508 33732 -4488
rect 33648 -4516 33668 -4508
rect 33676 -4516 33704 -4508
rect 33712 -4516 33732 -4508
rect 33768 -4508 33852 -4488
rect 33768 -4516 33788 -4508
rect 33796 -4516 33824 -4508
rect 33832 -4516 33852 -4508
rect 33888 -4508 33972 -4488
rect 33888 -4516 33908 -4508
rect 33916 -4516 33944 -4508
rect 33952 -4516 33972 -4508
rect 34008 -4508 34092 -4488
rect 34008 -4516 34028 -4508
rect 34036 -4516 34064 -4508
rect 34072 -4516 34092 -4508
rect 34128 -4508 34212 -4488
rect 34128 -4516 34148 -4508
rect 34156 -4516 34184 -4508
rect 34192 -4516 34212 -4508
rect 34248 -4508 34332 -4488
rect 34248 -4516 34268 -4508
rect 34276 -4516 34304 -4508
rect 34312 -4516 34332 -4508
rect 34368 -4508 34452 -4488
rect 34368 -4516 34388 -4508
rect 34396 -4516 34424 -4508
rect 34432 -4516 34452 -4508
rect 34488 -4508 34572 -4488
rect 34488 -4516 34508 -4508
rect 34516 -4516 34544 -4508
rect 34552 -4516 34572 -4508
rect 34608 -4508 34692 -4488
rect 34608 -4516 34628 -4508
rect 34636 -4516 34664 -4508
rect 34672 -4516 34692 -4508
rect 34728 -4508 34812 -4488
rect 34728 -4516 34748 -4508
rect 34756 -4516 34784 -4508
rect 34792 -4516 34812 -4508
rect 34848 -4508 34932 -4488
rect 34848 -4516 34868 -4508
rect 34876 -4516 34904 -4508
rect 34912 -4516 34932 -4508
rect 34968 -4508 35052 -4488
rect 34968 -4516 34988 -4508
rect 34996 -4516 35024 -4508
rect 35032 -4516 35052 -4508
rect 35088 -4508 35172 -4488
rect 35088 -4516 35108 -4508
rect 35116 -4516 35144 -4508
rect 35152 -4516 35172 -4508
rect 35208 -4508 35292 -4488
rect 35208 -4516 35228 -4508
rect 35236 -4516 35264 -4508
rect 35272 -4516 35292 -4508
rect 35328 -4508 35412 -4488
rect 35328 -4516 35348 -4508
rect 35356 -4516 35384 -4508
rect 35392 -4516 35412 -4508
rect 35448 -4508 35532 -4488
rect 35448 -4516 35468 -4508
rect 35476 -4516 35504 -4508
rect 35512 -4516 35532 -4508
rect 35568 -4508 35652 -4488
rect 35568 -4516 35588 -4508
rect 35596 -4516 35624 -4508
rect 35632 -4516 35652 -4508
rect 35688 -4508 35772 -4488
rect 35688 -4516 35708 -4508
rect 35716 -4516 35744 -4508
rect 35752 -4516 35772 -4508
rect 35808 -4508 35892 -4488
rect 35808 -4516 35828 -4508
rect 35836 -4516 35864 -4508
rect 35872 -4516 35892 -4508
rect 35928 -4508 36012 -4488
rect 35928 -4516 35948 -4508
rect 35956 -4516 35984 -4508
rect 35992 -4516 36012 -4508
rect 36048 -4508 36132 -4488
rect 36048 -4516 36068 -4508
rect 36076 -4516 36104 -4508
rect 36112 -4516 36132 -4508
rect 36168 -4508 36252 -4488
rect 36168 -4516 36188 -4508
rect 36196 -4516 36224 -4508
rect 36232 -4516 36252 -4508
rect 36288 -4508 36372 -4488
rect 36288 -4516 36308 -4508
rect 36316 -4516 36344 -4508
rect 36352 -4516 36372 -4508
rect 36408 -4508 36492 -4488
rect 36408 -4516 36428 -4508
rect 36436 -4516 36464 -4508
rect 36472 -4516 36492 -4508
rect 36528 -4508 36612 -4488
rect 36528 -4516 36548 -4508
rect 36556 -4516 36584 -4508
rect 36592 -4516 36612 -4508
rect 36648 -4508 36732 -4488
rect 36648 -4516 36668 -4508
rect 36676 -4516 36704 -4508
rect 36712 -4516 36732 -4508
rect 36768 -4508 36852 -4488
rect 36768 -4516 36788 -4508
rect 36796 -4516 36824 -4508
rect 36832 -4516 36852 -4508
rect 36888 -4508 36972 -4488
rect 36888 -4516 36908 -4508
rect 36916 -4516 36944 -4508
rect 36952 -4516 36972 -4508
rect 37008 -4508 37092 -4488
rect 37008 -4516 37028 -4508
rect 37036 -4516 37064 -4508
rect 37072 -4516 37092 -4508
rect 37128 -4508 37212 -4488
rect 37128 -4516 37148 -4508
rect 37156 -4516 37184 -4508
rect 37192 -4516 37212 -4508
rect 37248 -4508 37332 -4488
rect 37248 -4516 37268 -4508
rect 37276 -4516 37304 -4508
rect 37312 -4516 37332 -4508
rect 37368 -4508 37452 -4488
rect 37368 -4516 37388 -4508
rect 37396 -4516 37424 -4508
rect 37432 -4516 37452 -4508
rect 37488 -4508 37572 -4488
rect 37488 -4516 37508 -4508
rect 37516 -4516 37544 -4508
rect 37552 -4516 37572 -4508
rect 37608 -4508 37692 -4488
rect 37608 -4516 37628 -4508
rect 37636 -4516 37664 -4508
rect 37672 -4516 37692 -4508
rect 37728 -4508 37812 -4488
rect 37728 -4516 37748 -4508
rect 37756 -4516 37784 -4508
rect 37792 -4516 37812 -4508
rect 37848 -4508 37932 -4488
rect 37848 -4516 37868 -4508
rect 37876 -4516 37904 -4508
rect 37912 -4516 37932 -4508
rect 37968 -4508 38052 -4488
rect 37968 -4516 37988 -4508
rect 37996 -4516 38024 -4508
rect 38032 -4516 38052 -4508
rect 38088 -4508 38172 -4488
rect 38088 -4516 38108 -4508
rect 38116 -4516 38144 -4508
rect 38152 -4516 38172 -4508
rect 38208 -4508 38292 -4488
rect 38208 -4516 38228 -4508
rect 38236 -4516 38264 -4508
rect 38272 -4516 38292 -4508
rect 38328 -4508 38412 -4488
rect 38328 -4516 38348 -4508
rect 38356 -4516 38384 -4508
rect 38392 -4516 38412 -4508
rect 38448 -4508 38532 -4488
rect 38448 -4516 38468 -4508
rect 38476 -4516 38504 -4508
rect 38512 -4516 38532 -4508
rect 38568 -4508 38652 -4488
rect 38568 -4516 38588 -4508
rect 38596 -4516 38624 -4508
rect 38632 -4516 38652 -4508
rect 38688 -4508 38772 -4488
rect 38688 -4516 38708 -4508
rect 38716 -4516 38744 -4508
rect 38752 -4516 38772 -4508
rect 38808 -4508 38892 -4488
rect 38808 -4516 38828 -4508
rect 38836 -4516 38864 -4508
rect 38872 -4516 38892 -4508
rect 38928 -4508 39012 -4488
rect 38928 -4516 38948 -4508
rect 38956 -4516 38984 -4508
rect 38992 -4516 39012 -4508
rect 39048 -4508 39132 -4488
rect 39048 -4516 39068 -4508
rect 39076 -4516 39104 -4508
rect 39112 -4516 39132 -4508
rect 39168 -4508 39252 -4488
rect 39168 -4516 39188 -4508
rect 39196 -4516 39224 -4508
rect 39232 -4516 39252 -4508
rect 39288 -4508 39372 -4488
rect 39288 -4516 39308 -4508
rect 39316 -4516 39344 -4508
rect 39352 -4516 39372 -4508
rect 39408 -4508 39492 -4488
rect 39408 -4516 39428 -4508
rect 39436 -4516 39464 -4508
rect 39472 -4516 39492 -4508
rect 39528 -4508 39612 -4488
rect 39528 -4516 39548 -4508
rect 39556 -4516 39584 -4508
rect 39592 -4516 39612 -4508
rect 39648 -4508 39732 -4488
rect 39648 -4516 39668 -4508
rect 39676 -4516 39704 -4508
rect 39712 -4516 39732 -4508
rect 39768 -4508 39852 -4488
rect 39768 -4516 39788 -4508
rect 39796 -4516 39824 -4508
rect 39832 -4516 39852 -4508
rect 39888 -4508 39972 -4488
rect 39888 -4516 39908 -4508
rect 39916 -4516 39944 -4508
rect 39952 -4516 39972 -4508
rect 40008 -4508 40092 -4488
rect 40008 -4516 40028 -4508
rect 40036 -4516 40064 -4508
rect 40072 -4516 40092 -4508
rect 40128 -4508 40212 -4488
rect 40128 -4516 40148 -4508
rect 40156 -4516 40184 -4508
rect 40192 -4516 40212 -4508
rect 40248 -4508 40332 -4488
rect 40248 -4516 40268 -4508
rect 40276 -4516 40304 -4508
rect 40312 -4516 40332 -4508
rect 40368 -4508 40452 -4488
rect 40368 -4516 40388 -4508
rect 40396 -4516 40424 -4508
rect 40432 -4516 40452 -4508
rect 40488 -4508 40572 -4488
rect 40488 -4516 40508 -4508
rect 40516 -4516 40544 -4508
rect 40552 -4516 40572 -4508
rect 40608 -4508 40692 -4488
rect 40608 -4516 40628 -4508
rect 40636 -4516 40664 -4508
rect 40672 -4516 40692 -4508
rect 40728 -4508 40812 -4488
rect 40728 -4516 40748 -4508
rect 40756 -4516 40784 -4508
rect 40792 -4516 40812 -4508
rect 40848 -4508 40932 -4488
rect 40848 -4516 40868 -4508
rect 40876 -4516 40904 -4508
rect 40912 -4516 40932 -4508
rect 40968 -4508 41052 -4488
rect 40968 -4516 40988 -4508
rect 40996 -4516 41024 -4508
rect 41032 -4516 41052 -4508
rect 41088 -4508 41172 -4488
rect 41088 -4516 41108 -4508
rect 41116 -4516 41144 -4508
rect 41152 -4516 41172 -4508
rect 41208 -4508 41292 -4488
rect 41208 -4516 41228 -4508
rect 41236 -4516 41264 -4508
rect 41272 -4516 41292 -4508
rect 41328 -4508 41412 -4488
rect 41328 -4516 41348 -4508
rect 41356 -4516 41384 -4508
rect 41392 -4516 41412 -4508
rect 41448 -4508 41532 -4488
rect 41448 -4516 41468 -4508
rect 41476 -4516 41504 -4508
rect 41512 -4516 41532 -4508
rect 41568 -4508 41652 -4488
rect 41568 -4516 41588 -4508
rect 41596 -4516 41624 -4508
rect 41632 -4516 41652 -4508
rect 41688 -4508 41772 -4488
rect 41688 -4516 41708 -4508
rect 41716 -4516 41744 -4508
rect 41752 -4516 41772 -4508
rect 41808 -4508 41892 -4488
rect 41808 -4516 41828 -4508
rect 41836 -4516 41864 -4508
rect 41872 -4516 41892 -4508
rect 41928 -4508 42012 -4488
rect 41928 -4516 41948 -4508
rect 41956 -4516 41984 -4508
rect 41992 -4516 42012 -4508
rect 42048 -4508 42132 -4488
rect 42048 -4516 42068 -4508
rect 42076 -4516 42104 -4508
rect 42112 -4516 42132 -4508
rect 42168 -4508 42252 -4488
rect 42168 -4516 42188 -4508
rect 42196 -4516 42224 -4508
rect 42232 -4516 42252 -4508
rect 42288 -4508 42372 -4488
rect 42288 -4516 42308 -4508
rect 42316 -4516 42344 -4508
rect 42352 -4516 42372 -4508
rect 42408 -4508 42492 -4488
rect 42408 -4516 42428 -4508
rect 42436 -4516 42464 -4508
rect 42472 -4516 42492 -4508
rect 42528 -4508 42612 -4488
rect 42528 -4516 42548 -4508
rect 42556 -4516 42584 -4508
rect 42592 -4516 42612 -4508
rect 42648 -4508 42732 -4488
rect 42648 -4516 42668 -4508
rect 42676 -4516 42704 -4508
rect 42712 -4516 42732 -4508
rect 42768 -4508 42852 -4488
rect 42768 -4516 42788 -4508
rect 42796 -4516 42824 -4508
rect 42832 -4516 42852 -4508
rect 42888 -4508 42972 -4488
rect 42888 -4516 42908 -4508
rect 42916 -4516 42944 -4508
rect 42952 -4516 42972 -4508
rect 43008 -4508 43092 -4488
rect 43008 -4516 43028 -4508
rect 43036 -4516 43064 -4508
rect 43072 -4516 43092 -4508
rect 43128 -4508 43212 -4488
rect 43128 -4516 43148 -4508
rect 43156 -4516 43184 -4508
rect 43192 -4516 43212 -4508
rect 43248 -4508 43332 -4488
rect 43248 -4516 43268 -4508
rect 43276 -4516 43304 -4508
rect 43312 -4516 43332 -4508
rect 43368 -4508 43452 -4488
rect 43368 -4516 43388 -4508
rect 43396 -4516 43424 -4508
rect 43432 -4516 43452 -4508
rect 43488 -4508 43572 -4488
rect 43488 -4516 43508 -4508
rect 43516 -4516 43544 -4508
rect 43552 -4516 43572 -4508
rect 43608 -4508 43692 -4488
rect 43608 -4516 43628 -4508
rect 43636 -4516 43664 -4508
rect 43672 -4516 43692 -4508
rect 43728 -4508 43812 -4488
rect 43728 -4516 43748 -4508
rect 43756 -4516 43784 -4508
rect 43792 -4516 43812 -4508
rect 43848 -4508 43932 -4488
rect 43848 -4516 43868 -4508
rect 43876 -4516 43904 -4508
rect 43912 -4516 43932 -4508
rect 43968 -4508 44052 -4488
rect 43968 -4516 43988 -4508
rect 43996 -4516 44024 -4508
rect 44032 -4516 44052 -4508
rect 44088 -4508 44172 -4488
rect 44088 -4516 44108 -4508
rect 44116 -4516 44144 -4508
rect 44152 -4516 44172 -4508
rect 44208 -4508 44292 -4488
rect 44208 -4516 44228 -4508
rect 44236 -4516 44264 -4508
rect 44272 -4516 44292 -4508
rect 44328 -4508 44412 -4488
rect 44328 -4516 44348 -4508
rect 44356 -4516 44384 -4508
rect 44392 -4516 44412 -4508
rect 44448 -4508 44532 -4488
rect 44448 -4516 44468 -4508
rect 44476 -4516 44504 -4508
rect 44512 -4516 44532 -4508
rect 44568 -4508 44652 -4488
rect 44568 -4516 44588 -4508
rect 44596 -4516 44624 -4508
rect 44632 -4516 44652 -4508
rect 44688 -4508 44772 -4488
rect 44688 -4516 44708 -4508
rect 44716 -4516 44744 -4508
rect 44752 -4516 44772 -4508
rect 44808 -4508 44892 -4488
rect 44808 -4516 44828 -4508
rect 44836 -4516 44864 -4508
rect 44872 -4516 44892 -4508
rect 44928 -4508 45012 -4488
rect 44928 -4516 44948 -4508
rect 44956 -4516 44984 -4508
rect 44992 -4516 45012 -4508
rect 45048 -4508 45132 -4488
rect 45048 -4516 45068 -4508
rect 45076 -4516 45104 -4508
rect 45112 -4516 45132 -4508
rect 45168 -4508 45252 -4488
rect 45168 -4516 45188 -4508
rect 45196 -4516 45224 -4508
rect 45232 -4516 45252 -4508
rect 45288 -4508 45372 -4488
rect 45288 -4516 45308 -4508
rect 45316 -4516 45344 -4508
rect 45352 -4516 45372 -4508
rect 45408 -4508 45492 -4488
rect 45408 -4516 45428 -4508
rect 45436 -4516 45464 -4508
rect 45472 -4516 45492 -4508
rect 45528 -4508 45612 -4488
rect 45528 -4516 45548 -4508
rect 45556 -4516 45584 -4508
rect 45592 -4516 45612 -4508
rect 25876 -4544 25932 -4516
rect 25996 -4544 26052 -4516
rect 26116 -4544 26172 -4516
rect 26236 -4544 26292 -4516
rect 26356 -4544 26412 -4516
rect 26476 -4544 26532 -4516
rect 26596 -4544 26652 -4516
rect 26716 -4544 26772 -4516
rect 26836 -4544 26892 -4516
rect 26956 -4544 27012 -4516
rect 27076 -4544 27132 -4516
rect 27196 -4544 27252 -4516
rect 27316 -4544 27372 -4516
rect 27436 -4544 27492 -4516
rect 27556 -4544 27612 -4516
rect 27676 -4544 27732 -4516
rect 27796 -4544 27852 -4516
rect 27916 -4544 27972 -4516
rect 28036 -4544 28092 -4516
rect 28156 -4544 28212 -4516
rect 28276 -4544 28332 -4516
rect 28396 -4544 28452 -4516
rect 28516 -4544 28572 -4516
rect 28636 -4544 28692 -4516
rect 28756 -4544 28812 -4516
rect 28876 -4544 28932 -4516
rect 28996 -4544 29052 -4516
rect 29116 -4544 29172 -4516
rect 29236 -4544 29292 -4516
rect 29356 -4544 29412 -4516
rect 29476 -4544 29532 -4516
rect 29596 -4544 29652 -4516
rect 29716 -4544 29772 -4516
rect 29836 -4544 29892 -4516
rect 29956 -4544 30012 -4516
rect 30076 -4544 30132 -4516
rect 30196 -4544 30252 -4516
rect 30316 -4544 30372 -4516
rect 30436 -4544 30492 -4516
rect 30556 -4544 30612 -4516
rect 30676 -4544 30732 -4516
rect 30796 -4544 30852 -4516
rect 30916 -4544 30972 -4516
rect 31036 -4544 31092 -4516
rect 31156 -4544 31212 -4516
rect 31276 -4544 31332 -4516
rect 31396 -4544 31452 -4516
rect 31516 -4544 31572 -4516
rect 31636 -4544 31692 -4516
rect 31756 -4544 31812 -4516
rect 31876 -4544 31932 -4516
rect 31996 -4544 32052 -4516
rect 32116 -4544 32172 -4516
rect 32236 -4544 32292 -4516
rect 32356 -4544 32412 -4516
rect 32476 -4544 32532 -4516
rect 32596 -4544 32652 -4516
rect 32716 -4544 32772 -4516
rect 32836 -4544 32892 -4516
rect 32956 -4544 33012 -4516
rect 33076 -4544 33132 -4516
rect 33196 -4544 33252 -4516
rect 33316 -4544 33372 -4516
rect 33436 -4544 33492 -4516
rect 33556 -4544 33612 -4516
rect 33676 -4544 33732 -4516
rect 33796 -4544 33852 -4516
rect 33916 -4544 33972 -4516
rect 34036 -4544 34092 -4516
rect 34156 -4544 34212 -4516
rect 34276 -4544 34332 -4516
rect 34396 -4544 34452 -4516
rect 34516 -4544 34572 -4516
rect 34636 -4544 34692 -4516
rect 34756 -4544 34812 -4516
rect 34876 -4544 34932 -4516
rect 34996 -4544 35052 -4516
rect 35116 -4544 35172 -4516
rect 35236 -4544 35292 -4516
rect 35356 -4544 35412 -4516
rect 35476 -4544 35532 -4516
rect 35596 -4544 35652 -4516
rect 35716 -4544 35772 -4516
rect 35836 -4544 35892 -4516
rect 35956 -4544 36012 -4516
rect 36076 -4544 36132 -4516
rect 36196 -4544 36252 -4516
rect 36316 -4544 36372 -4516
rect 36436 -4544 36492 -4516
rect 36556 -4544 36612 -4516
rect 36676 -4544 36732 -4516
rect 36796 -4544 36852 -4516
rect 36916 -4544 36972 -4516
rect 37036 -4544 37092 -4516
rect 37156 -4544 37212 -4516
rect 37276 -4544 37332 -4516
rect 37396 -4544 37452 -4516
rect 37516 -4544 37572 -4516
rect 37636 -4544 37692 -4516
rect 37756 -4544 37812 -4516
rect 37876 -4544 37932 -4516
rect 37996 -4544 38052 -4516
rect 38116 -4544 38172 -4516
rect 38236 -4544 38292 -4516
rect 38356 -4544 38412 -4516
rect 38476 -4544 38532 -4516
rect 38596 -4544 38652 -4516
rect 38716 -4544 38772 -4516
rect 38836 -4544 38892 -4516
rect 38956 -4544 39012 -4516
rect 39076 -4544 39132 -4516
rect 39196 -4544 39252 -4516
rect 39316 -4544 39372 -4516
rect 39436 -4544 39492 -4516
rect 39556 -4544 39612 -4516
rect 39676 -4544 39732 -4516
rect 39796 -4544 39852 -4516
rect 39916 -4544 39972 -4516
rect 40036 -4544 40092 -4516
rect 40156 -4544 40212 -4516
rect 40276 -4544 40332 -4516
rect 40396 -4544 40452 -4516
rect 40516 -4544 40572 -4516
rect 40636 -4544 40692 -4516
rect 40756 -4544 40812 -4516
rect 40876 -4544 40932 -4516
rect 40996 -4544 41052 -4516
rect 41116 -4544 41172 -4516
rect 41236 -4544 41292 -4516
rect 41356 -4544 41412 -4516
rect 41476 -4544 41532 -4516
rect 41596 -4544 41652 -4516
rect 41716 -4544 41772 -4516
rect 41836 -4544 41892 -4516
rect 41956 -4544 42012 -4516
rect 42076 -4544 42132 -4516
rect 42196 -4544 42252 -4516
rect 42316 -4544 42372 -4516
rect 42436 -4544 42492 -4516
rect 42556 -4544 42612 -4516
rect 42676 -4544 42732 -4516
rect 42796 -4544 42852 -4516
rect 42916 -4544 42972 -4516
rect 43036 -4544 43092 -4516
rect 43156 -4544 43212 -4516
rect 43276 -4544 43332 -4516
rect 43396 -4544 43452 -4516
rect 43516 -4544 43572 -4516
rect 43636 -4544 43692 -4516
rect 43756 -4544 43812 -4516
rect 43876 -4544 43932 -4516
rect 43996 -4544 44052 -4516
rect 44116 -4544 44172 -4516
rect 44236 -4544 44292 -4516
rect 44356 -4544 44412 -4516
rect 44476 -4544 44532 -4516
rect 44596 -4544 44652 -4516
rect 44716 -4544 44772 -4516
rect 44836 -4544 44892 -4516
rect 44956 -4544 45012 -4516
rect 45076 -4544 45132 -4516
rect 45196 -4544 45252 -4516
rect 45316 -4544 45372 -4516
rect 45436 -4544 45492 -4516
rect 45556 -4544 45612 -4516
rect 25848 -4688 25932 -4668
rect 25848 -4696 25868 -4688
rect 25876 -4696 25904 -4688
rect 25912 -4696 25932 -4688
rect 25968 -4688 26052 -4668
rect 25968 -4696 25988 -4688
rect 25996 -4696 26024 -4688
rect 26032 -4696 26052 -4688
rect 26088 -4688 26172 -4668
rect 26088 -4696 26108 -4688
rect 26116 -4696 26144 -4688
rect 26152 -4696 26172 -4688
rect 26208 -4688 26292 -4668
rect 26208 -4696 26228 -4688
rect 26236 -4696 26264 -4688
rect 26272 -4696 26292 -4688
rect 26328 -4688 26412 -4668
rect 26328 -4696 26348 -4688
rect 26356 -4696 26384 -4688
rect 26392 -4696 26412 -4688
rect 26448 -4688 26532 -4668
rect 26448 -4696 26468 -4688
rect 26476 -4696 26504 -4688
rect 26512 -4696 26532 -4688
rect 26568 -4688 26652 -4668
rect 26568 -4696 26588 -4688
rect 26596 -4696 26624 -4688
rect 26632 -4696 26652 -4688
rect 26688 -4688 26772 -4668
rect 26688 -4696 26708 -4688
rect 26716 -4696 26744 -4688
rect 26752 -4696 26772 -4688
rect 26808 -4688 26892 -4668
rect 26808 -4696 26828 -4688
rect 26836 -4696 26864 -4688
rect 26872 -4696 26892 -4688
rect 26928 -4688 27012 -4668
rect 26928 -4696 26948 -4688
rect 26956 -4696 26984 -4688
rect 26992 -4696 27012 -4688
rect 27048 -4688 27132 -4668
rect 27048 -4696 27068 -4688
rect 27076 -4696 27104 -4688
rect 27112 -4696 27132 -4688
rect 27168 -4688 27252 -4668
rect 27168 -4696 27188 -4688
rect 27196 -4696 27224 -4688
rect 27232 -4696 27252 -4688
rect 27288 -4688 27372 -4668
rect 27288 -4696 27308 -4688
rect 27316 -4696 27344 -4688
rect 27352 -4696 27372 -4688
rect 27408 -4688 27492 -4668
rect 27408 -4696 27428 -4688
rect 27436 -4696 27464 -4688
rect 27472 -4696 27492 -4688
rect 27528 -4688 27612 -4668
rect 27528 -4696 27548 -4688
rect 27556 -4696 27584 -4688
rect 27592 -4696 27612 -4688
rect 27648 -4688 27732 -4668
rect 27648 -4696 27668 -4688
rect 27676 -4696 27704 -4688
rect 27712 -4696 27732 -4688
rect 27768 -4688 27852 -4668
rect 27768 -4696 27788 -4688
rect 27796 -4696 27824 -4688
rect 27832 -4696 27852 -4688
rect 27888 -4688 27972 -4668
rect 27888 -4696 27908 -4688
rect 27916 -4696 27944 -4688
rect 27952 -4696 27972 -4688
rect 28008 -4688 28092 -4668
rect 28008 -4696 28028 -4688
rect 28036 -4696 28064 -4688
rect 28072 -4696 28092 -4688
rect 28128 -4688 28212 -4668
rect 28128 -4696 28148 -4688
rect 28156 -4696 28184 -4688
rect 28192 -4696 28212 -4688
rect 28248 -4688 28332 -4668
rect 28248 -4696 28268 -4688
rect 28276 -4696 28304 -4688
rect 28312 -4696 28332 -4688
rect 28368 -4688 28452 -4668
rect 28368 -4696 28388 -4688
rect 28396 -4696 28424 -4688
rect 28432 -4696 28452 -4688
rect 28488 -4688 28572 -4668
rect 28488 -4696 28508 -4688
rect 28516 -4696 28544 -4688
rect 28552 -4696 28572 -4688
rect 28608 -4688 28692 -4668
rect 28608 -4696 28628 -4688
rect 28636 -4696 28664 -4688
rect 28672 -4696 28692 -4688
rect 28728 -4688 28812 -4668
rect 28728 -4696 28748 -4688
rect 28756 -4696 28784 -4688
rect 28792 -4696 28812 -4688
rect 28848 -4688 28932 -4668
rect 28848 -4696 28868 -4688
rect 28876 -4696 28904 -4688
rect 28912 -4696 28932 -4688
rect 28968 -4688 29052 -4668
rect 28968 -4696 28988 -4688
rect 28996 -4696 29024 -4688
rect 29032 -4696 29052 -4688
rect 29088 -4688 29172 -4668
rect 29088 -4696 29108 -4688
rect 29116 -4696 29144 -4688
rect 29152 -4696 29172 -4688
rect 29208 -4688 29292 -4668
rect 29208 -4696 29228 -4688
rect 29236 -4696 29264 -4688
rect 29272 -4696 29292 -4688
rect 29328 -4688 29412 -4668
rect 29328 -4696 29348 -4688
rect 29356 -4696 29384 -4688
rect 29392 -4696 29412 -4688
rect 29448 -4688 29532 -4668
rect 29448 -4696 29468 -4688
rect 29476 -4696 29504 -4688
rect 29512 -4696 29532 -4688
rect 29568 -4688 29652 -4668
rect 29568 -4696 29588 -4688
rect 29596 -4696 29624 -4688
rect 29632 -4696 29652 -4688
rect 29688 -4688 29772 -4668
rect 29688 -4696 29708 -4688
rect 29716 -4696 29744 -4688
rect 29752 -4696 29772 -4688
rect 29808 -4688 29892 -4668
rect 29808 -4696 29828 -4688
rect 29836 -4696 29864 -4688
rect 29872 -4696 29892 -4688
rect 29928 -4688 30012 -4668
rect 29928 -4696 29948 -4688
rect 29956 -4696 29984 -4688
rect 29992 -4696 30012 -4688
rect 30048 -4688 30132 -4668
rect 30048 -4696 30068 -4688
rect 30076 -4696 30104 -4688
rect 30112 -4696 30132 -4688
rect 30168 -4688 30252 -4668
rect 30168 -4696 30188 -4688
rect 30196 -4696 30224 -4688
rect 30232 -4696 30252 -4688
rect 30288 -4688 30372 -4668
rect 30288 -4696 30308 -4688
rect 30316 -4696 30344 -4688
rect 30352 -4696 30372 -4688
rect 30408 -4688 30492 -4668
rect 30408 -4696 30428 -4688
rect 30436 -4696 30464 -4688
rect 30472 -4696 30492 -4688
rect 30528 -4688 30612 -4668
rect 30528 -4696 30548 -4688
rect 30556 -4696 30584 -4688
rect 30592 -4696 30612 -4688
rect 30648 -4688 30732 -4668
rect 30648 -4696 30668 -4688
rect 30676 -4696 30704 -4688
rect 30712 -4696 30732 -4688
rect 30768 -4688 30852 -4668
rect 30768 -4696 30788 -4688
rect 30796 -4696 30824 -4688
rect 30832 -4696 30852 -4688
rect 30888 -4688 30972 -4668
rect 30888 -4696 30908 -4688
rect 30916 -4696 30944 -4688
rect 30952 -4696 30972 -4688
rect 31008 -4688 31092 -4668
rect 31008 -4696 31028 -4688
rect 31036 -4696 31064 -4688
rect 31072 -4696 31092 -4688
rect 31128 -4688 31212 -4668
rect 31128 -4696 31148 -4688
rect 31156 -4696 31184 -4688
rect 31192 -4696 31212 -4688
rect 31248 -4688 31332 -4668
rect 31248 -4696 31268 -4688
rect 31276 -4696 31304 -4688
rect 31312 -4696 31332 -4688
rect 31368 -4688 31452 -4668
rect 31368 -4696 31388 -4688
rect 31396 -4696 31424 -4688
rect 31432 -4696 31452 -4688
rect 31488 -4688 31572 -4668
rect 31488 -4696 31508 -4688
rect 31516 -4696 31544 -4688
rect 31552 -4696 31572 -4688
rect 31608 -4688 31692 -4668
rect 31608 -4696 31628 -4688
rect 31636 -4696 31664 -4688
rect 31672 -4696 31692 -4688
rect 31728 -4688 31812 -4668
rect 31728 -4696 31748 -4688
rect 31756 -4696 31784 -4688
rect 31792 -4696 31812 -4688
rect 31848 -4688 31932 -4668
rect 31848 -4696 31868 -4688
rect 31876 -4696 31904 -4688
rect 31912 -4696 31932 -4688
rect 31968 -4688 32052 -4668
rect 31968 -4696 31988 -4688
rect 31996 -4696 32024 -4688
rect 32032 -4696 32052 -4688
rect 32088 -4688 32172 -4668
rect 32088 -4696 32108 -4688
rect 32116 -4696 32144 -4688
rect 32152 -4696 32172 -4688
rect 32208 -4688 32292 -4668
rect 32208 -4696 32228 -4688
rect 32236 -4696 32264 -4688
rect 32272 -4696 32292 -4688
rect 32328 -4688 32412 -4668
rect 32328 -4696 32348 -4688
rect 32356 -4696 32384 -4688
rect 32392 -4696 32412 -4688
rect 32448 -4688 32532 -4668
rect 32448 -4696 32468 -4688
rect 32476 -4696 32504 -4688
rect 32512 -4696 32532 -4688
rect 32568 -4688 32652 -4668
rect 32568 -4696 32588 -4688
rect 32596 -4696 32624 -4688
rect 32632 -4696 32652 -4688
rect 32688 -4688 32772 -4668
rect 32688 -4696 32708 -4688
rect 32716 -4696 32744 -4688
rect 32752 -4696 32772 -4688
rect 32808 -4688 32892 -4668
rect 32808 -4696 32828 -4688
rect 32836 -4696 32864 -4688
rect 32872 -4696 32892 -4688
rect 32928 -4688 33012 -4668
rect 32928 -4696 32948 -4688
rect 32956 -4696 32984 -4688
rect 32992 -4696 33012 -4688
rect 33048 -4688 33132 -4668
rect 33048 -4696 33068 -4688
rect 33076 -4696 33104 -4688
rect 33112 -4696 33132 -4688
rect 33168 -4688 33252 -4668
rect 33168 -4696 33188 -4688
rect 33196 -4696 33224 -4688
rect 33232 -4696 33252 -4688
rect 33288 -4688 33372 -4668
rect 33288 -4696 33308 -4688
rect 33316 -4696 33344 -4688
rect 33352 -4696 33372 -4688
rect 33408 -4688 33492 -4668
rect 33408 -4696 33428 -4688
rect 33436 -4696 33464 -4688
rect 33472 -4696 33492 -4688
rect 33528 -4688 33612 -4668
rect 33528 -4696 33548 -4688
rect 33556 -4696 33584 -4688
rect 33592 -4696 33612 -4688
rect 33648 -4688 33732 -4668
rect 33648 -4696 33668 -4688
rect 33676 -4696 33704 -4688
rect 33712 -4696 33732 -4688
rect 33768 -4688 33852 -4668
rect 33768 -4696 33788 -4688
rect 33796 -4696 33824 -4688
rect 33832 -4696 33852 -4688
rect 33888 -4688 33972 -4668
rect 33888 -4696 33908 -4688
rect 33916 -4696 33944 -4688
rect 33952 -4696 33972 -4688
rect 34008 -4688 34092 -4668
rect 34008 -4696 34028 -4688
rect 34036 -4696 34064 -4688
rect 34072 -4696 34092 -4688
rect 34128 -4688 34212 -4668
rect 34128 -4696 34148 -4688
rect 34156 -4696 34184 -4688
rect 34192 -4696 34212 -4688
rect 34248 -4688 34332 -4668
rect 34248 -4696 34268 -4688
rect 34276 -4696 34304 -4688
rect 34312 -4696 34332 -4688
rect 34368 -4688 34452 -4668
rect 34368 -4696 34388 -4688
rect 34396 -4696 34424 -4688
rect 34432 -4696 34452 -4688
rect 34488 -4688 34572 -4668
rect 34488 -4696 34508 -4688
rect 34516 -4696 34544 -4688
rect 34552 -4696 34572 -4688
rect 34608 -4688 34692 -4668
rect 34608 -4696 34628 -4688
rect 34636 -4696 34664 -4688
rect 34672 -4696 34692 -4688
rect 34728 -4688 34812 -4668
rect 34728 -4696 34748 -4688
rect 34756 -4696 34784 -4688
rect 34792 -4696 34812 -4688
rect 34848 -4688 34932 -4668
rect 34848 -4696 34868 -4688
rect 34876 -4696 34904 -4688
rect 34912 -4696 34932 -4688
rect 34968 -4688 35052 -4668
rect 34968 -4696 34988 -4688
rect 34996 -4696 35024 -4688
rect 35032 -4696 35052 -4688
rect 35088 -4688 35172 -4668
rect 35088 -4696 35108 -4688
rect 35116 -4696 35144 -4688
rect 35152 -4696 35172 -4688
rect 35208 -4688 35292 -4668
rect 35208 -4696 35228 -4688
rect 35236 -4696 35264 -4688
rect 35272 -4696 35292 -4688
rect 35328 -4688 35412 -4668
rect 35328 -4696 35348 -4688
rect 35356 -4696 35384 -4688
rect 35392 -4696 35412 -4688
rect 35448 -4688 35532 -4668
rect 35448 -4696 35468 -4688
rect 35476 -4696 35504 -4688
rect 35512 -4696 35532 -4688
rect 35568 -4688 35652 -4668
rect 35568 -4696 35588 -4688
rect 35596 -4696 35624 -4688
rect 35632 -4696 35652 -4688
rect 35688 -4688 35772 -4668
rect 35688 -4696 35708 -4688
rect 35716 -4696 35744 -4688
rect 35752 -4696 35772 -4688
rect 35808 -4688 35892 -4668
rect 35808 -4696 35828 -4688
rect 35836 -4696 35864 -4688
rect 35872 -4696 35892 -4688
rect 35928 -4688 36012 -4668
rect 35928 -4696 35948 -4688
rect 35956 -4696 35984 -4688
rect 35992 -4696 36012 -4688
rect 36048 -4688 36132 -4668
rect 36048 -4696 36068 -4688
rect 36076 -4696 36104 -4688
rect 36112 -4696 36132 -4688
rect 36168 -4688 36252 -4668
rect 36168 -4696 36188 -4688
rect 36196 -4696 36224 -4688
rect 36232 -4696 36252 -4688
rect 36288 -4688 36372 -4668
rect 36288 -4696 36308 -4688
rect 36316 -4696 36344 -4688
rect 36352 -4696 36372 -4688
rect 36408 -4688 36492 -4668
rect 36408 -4696 36428 -4688
rect 36436 -4696 36464 -4688
rect 36472 -4696 36492 -4688
rect 36528 -4688 36612 -4668
rect 36528 -4696 36548 -4688
rect 36556 -4696 36584 -4688
rect 36592 -4696 36612 -4688
rect 36648 -4688 36732 -4668
rect 36648 -4696 36668 -4688
rect 36676 -4696 36704 -4688
rect 36712 -4696 36732 -4688
rect 36768 -4688 36852 -4668
rect 36768 -4696 36788 -4688
rect 36796 -4696 36824 -4688
rect 36832 -4696 36852 -4688
rect 36888 -4688 36972 -4668
rect 36888 -4696 36908 -4688
rect 36916 -4696 36944 -4688
rect 36952 -4696 36972 -4688
rect 37008 -4688 37092 -4668
rect 37008 -4696 37028 -4688
rect 37036 -4696 37064 -4688
rect 37072 -4696 37092 -4688
rect 37128 -4688 37212 -4668
rect 37128 -4696 37148 -4688
rect 37156 -4696 37184 -4688
rect 37192 -4696 37212 -4688
rect 37248 -4688 37332 -4668
rect 37248 -4696 37268 -4688
rect 37276 -4696 37304 -4688
rect 37312 -4696 37332 -4688
rect 37368 -4688 37452 -4668
rect 37368 -4696 37388 -4688
rect 37396 -4696 37424 -4688
rect 37432 -4696 37452 -4688
rect 37488 -4688 37572 -4668
rect 37488 -4696 37508 -4688
rect 37516 -4696 37544 -4688
rect 37552 -4696 37572 -4688
rect 37608 -4688 37692 -4668
rect 37608 -4696 37628 -4688
rect 37636 -4696 37664 -4688
rect 37672 -4696 37692 -4688
rect 37728 -4688 37812 -4668
rect 37728 -4696 37748 -4688
rect 37756 -4696 37784 -4688
rect 37792 -4696 37812 -4688
rect 37848 -4688 37932 -4668
rect 37848 -4696 37868 -4688
rect 37876 -4696 37904 -4688
rect 37912 -4696 37932 -4688
rect 37968 -4688 38052 -4668
rect 37968 -4696 37988 -4688
rect 37996 -4696 38024 -4688
rect 38032 -4696 38052 -4688
rect 38088 -4688 38172 -4668
rect 38088 -4696 38108 -4688
rect 38116 -4696 38144 -4688
rect 38152 -4696 38172 -4688
rect 38208 -4688 38292 -4668
rect 38208 -4696 38228 -4688
rect 38236 -4696 38264 -4688
rect 38272 -4696 38292 -4688
rect 38328 -4688 38412 -4668
rect 38328 -4696 38348 -4688
rect 38356 -4696 38384 -4688
rect 38392 -4696 38412 -4688
rect 38448 -4688 38532 -4668
rect 38448 -4696 38468 -4688
rect 38476 -4696 38504 -4688
rect 38512 -4696 38532 -4688
rect 38568 -4688 38652 -4668
rect 38568 -4696 38588 -4688
rect 38596 -4696 38624 -4688
rect 38632 -4696 38652 -4688
rect 38688 -4688 38772 -4668
rect 38688 -4696 38708 -4688
rect 38716 -4696 38744 -4688
rect 38752 -4696 38772 -4688
rect 38808 -4688 38892 -4668
rect 38808 -4696 38828 -4688
rect 38836 -4696 38864 -4688
rect 38872 -4696 38892 -4688
rect 38928 -4688 39012 -4668
rect 38928 -4696 38948 -4688
rect 38956 -4696 38984 -4688
rect 38992 -4696 39012 -4688
rect 39048 -4688 39132 -4668
rect 39048 -4696 39068 -4688
rect 39076 -4696 39104 -4688
rect 39112 -4696 39132 -4688
rect 39168 -4688 39252 -4668
rect 39168 -4696 39188 -4688
rect 39196 -4696 39224 -4688
rect 39232 -4696 39252 -4688
rect 39288 -4688 39372 -4668
rect 39288 -4696 39308 -4688
rect 39316 -4696 39344 -4688
rect 39352 -4696 39372 -4688
rect 39408 -4688 39492 -4668
rect 39408 -4696 39428 -4688
rect 39436 -4696 39464 -4688
rect 39472 -4696 39492 -4688
rect 39528 -4688 39612 -4668
rect 39528 -4696 39548 -4688
rect 39556 -4696 39584 -4688
rect 39592 -4696 39612 -4688
rect 39648 -4688 39732 -4668
rect 39648 -4696 39668 -4688
rect 39676 -4696 39704 -4688
rect 39712 -4696 39732 -4688
rect 39768 -4688 39852 -4668
rect 39768 -4696 39788 -4688
rect 39796 -4696 39824 -4688
rect 39832 -4696 39852 -4688
rect 39888 -4688 39972 -4668
rect 39888 -4696 39908 -4688
rect 39916 -4696 39944 -4688
rect 39952 -4696 39972 -4688
rect 40008 -4688 40092 -4668
rect 40008 -4696 40028 -4688
rect 40036 -4696 40064 -4688
rect 40072 -4696 40092 -4688
rect 40128 -4688 40212 -4668
rect 40128 -4696 40148 -4688
rect 40156 -4696 40184 -4688
rect 40192 -4696 40212 -4688
rect 40248 -4688 40332 -4668
rect 40248 -4696 40268 -4688
rect 40276 -4696 40304 -4688
rect 40312 -4696 40332 -4688
rect 40368 -4688 40452 -4668
rect 40368 -4696 40388 -4688
rect 40396 -4696 40424 -4688
rect 40432 -4696 40452 -4688
rect 40488 -4688 40572 -4668
rect 40488 -4696 40508 -4688
rect 40516 -4696 40544 -4688
rect 40552 -4696 40572 -4688
rect 40608 -4688 40692 -4668
rect 40608 -4696 40628 -4688
rect 40636 -4696 40664 -4688
rect 40672 -4696 40692 -4688
rect 40728 -4688 40812 -4668
rect 40728 -4696 40748 -4688
rect 40756 -4696 40784 -4688
rect 40792 -4696 40812 -4688
rect 40848 -4688 40932 -4668
rect 40848 -4696 40868 -4688
rect 40876 -4696 40904 -4688
rect 40912 -4696 40932 -4688
rect 40968 -4688 41052 -4668
rect 40968 -4696 40988 -4688
rect 40996 -4696 41024 -4688
rect 41032 -4696 41052 -4688
rect 41088 -4688 41172 -4668
rect 41088 -4696 41108 -4688
rect 41116 -4696 41144 -4688
rect 41152 -4696 41172 -4688
rect 41208 -4688 41292 -4668
rect 41208 -4696 41228 -4688
rect 41236 -4696 41264 -4688
rect 41272 -4696 41292 -4688
rect 41328 -4688 41412 -4668
rect 41328 -4696 41348 -4688
rect 41356 -4696 41384 -4688
rect 41392 -4696 41412 -4688
rect 41448 -4688 41532 -4668
rect 41448 -4696 41468 -4688
rect 41476 -4696 41504 -4688
rect 41512 -4696 41532 -4688
rect 41568 -4688 41652 -4668
rect 41568 -4696 41588 -4688
rect 41596 -4696 41624 -4688
rect 41632 -4696 41652 -4688
rect 41688 -4688 41772 -4668
rect 41688 -4696 41708 -4688
rect 41716 -4696 41744 -4688
rect 41752 -4696 41772 -4688
rect 41808 -4688 41892 -4668
rect 41808 -4696 41828 -4688
rect 41836 -4696 41864 -4688
rect 41872 -4696 41892 -4688
rect 41928 -4688 42012 -4668
rect 41928 -4696 41948 -4688
rect 41956 -4696 41984 -4688
rect 41992 -4696 42012 -4688
rect 42048 -4688 42132 -4668
rect 42048 -4696 42068 -4688
rect 42076 -4696 42104 -4688
rect 42112 -4696 42132 -4688
rect 42168 -4688 42252 -4668
rect 42168 -4696 42188 -4688
rect 42196 -4696 42224 -4688
rect 42232 -4696 42252 -4688
rect 42288 -4688 42372 -4668
rect 42288 -4696 42308 -4688
rect 42316 -4696 42344 -4688
rect 42352 -4696 42372 -4688
rect 42408 -4688 42492 -4668
rect 42408 -4696 42428 -4688
rect 42436 -4696 42464 -4688
rect 42472 -4696 42492 -4688
rect 42528 -4688 42612 -4668
rect 42528 -4696 42548 -4688
rect 42556 -4696 42584 -4688
rect 42592 -4696 42612 -4688
rect 42648 -4688 42732 -4668
rect 42648 -4696 42668 -4688
rect 42676 -4696 42704 -4688
rect 42712 -4696 42732 -4688
rect 42768 -4688 42852 -4668
rect 42768 -4696 42788 -4688
rect 42796 -4696 42824 -4688
rect 42832 -4696 42852 -4688
rect 42888 -4688 42972 -4668
rect 42888 -4696 42908 -4688
rect 42916 -4696 42944 -4688
rect 42952 -4696 42972 -4688
rect 43008 -4688 43092 -4668
rect 43008 -4696 43028 -4688
rect 43036 -4696 43064 -4688
rect 43072 -4696 43092 -4688
rect 43128 -4688 43212 -4668
rect 43128 -4696 43148 -4688
rect 43156 -4696 43184 -4688
rect 43192 -4696 43212 -4688
rect 43248 -4688 43332 -4668
rect 43248 -4696 43268 -4688
rect 43276 -4696 43304 -4688
rect 43312 -4696 43332 -4688
rect 43368 -4688 43452 -4668
rect 43368 -4696 43388 -4688
rect 43396 -4696 43424 -4688
rect 43432 -4696 43452 -4688
rect 43488 -4688 43572 -4668
rect 43488 -4696 43508 -4688
rect 43516 -4696 43544 -4688
rect 43552 -4696 43572 -4688
rect 43608 -4688 43692 -4668
rect 43608 -4696 43628 -4688
rect 43636 -4696 43664 -4688
rect 43672 -4696 43692 -4688
rect 43728 -4688 43812 -4668
rect 43728 -4696 43748 -4688
rect 43756 -4696 43784 -4688
rect 43792 -4696 43812 -4688
rect 43848 -4688 43932 -4668
rect 43848 -4696 43868 -4688
rect 43876 -4696 43904 -4688
rect 43912 -4696 43932 -4688
rect 43968 -4688 44052 -4668
rect 43968 -4696 43988 -4688
rect 43996 -4696 44024 -4688
rect 44032 -4696 44052 -4688
rect 44088 -4688 44172 -4668
rect 44088 -4696 44108 -4688
rect 44116 -4696 44144 -4688
rect 44152 -4696 44172 -4688
rect 44208 -4688 44292 -4668
rect 44208 -4696 44228 -4688
rect 44236 -4696 44264 -4688
rect 44272 -4696 44292 -4688
rect 44328 -4688 44412 -4668
rect 44328 -4696 44348 -4688
rect 44356 -4696 44384 -4688
rect 44392 -4696 44412 -4688
rect 44448 -4688 44532 -4668
rect 44448 -4696 44468 -4688
rect 44476 -4696 44504 -4688
rect 44512 -4696 44532 -4688
rect 44568 -4688 44652 -4668
rect 44568 -4696 44588 -4688
rect 44596 -4696 44624 -4688
rect 44632 -4696 44652 -4688
rect 44688 -4688 44772 -4668
rect 44688 -4696 44708 -4688
rect 44716 -4696 44744 -4688
rect 44752 -4696 44772 -4688
rect 44808 -4688 44892 -4668
rect 44808 -4696 44828 -4688
rect 44836 -4696 44864 -4688
rect 44872 -4696 44892 -4688
rect 44928 -4688 45012 -4668
rect 44928 -4696 44948 -4688
rect 44956 -4696 44984 -4688
rect 44992 -4696 45012 -4688
rect 45048 -4688 45132 -4668
rect 45048 -4696 45068 -4688
rect 45076 -4696 45104 -4688
rect 45112 -4696 45132 -4688
rect 45168 -4688 45252 -4668
rect 45168 -4696 45188 -4688
rect 45196 -4696 45224 -4688
rect 45232 -4696 45252 -4688
rect 45288 -4688 45372 -4668
rect 45288 -4696 45308 -4688
rect 45316 -4696 45344 -4688
rect 45352 -4696 45372 -4688
rect 45408 -4688 45492 -4668
rect 45408 -4696 45428 -4688
rect 45436 -4696 45464 -4688
rect 45472 -4696 45492 -4688
rect 45528 -4688 45612 -4668
rect 45528 -4696 45548 -4688
rect 45556 -4696 45584 -4688
rect 45592 -4696 45612 -4688
rect 25876 -4724 25932 -4696
rect 25996 -4724 26052 -4696
rect 26116 -4724 26172 -4696
rect 26236 -4724 26292 -4696
rect 26356 -4724 26412 -4696
rect 26476 -4724 26532 -4696
rect 26596 -4724 26652 -4696
rect 26716 -4724 26772 -4696
rect 26836 -4724 26892 -4696
rect 26956 -4724 27012 -4696
rect 27076 -4724 27132 -4696
rect 27196 -4724 27252 -4696
rect 27316 -4724 27372 -4696
rect 27436 -4724 27492 -4696
rect 27556 -4724 27612 -4696
rect 27676 -4724 27732 -4696
rect 27796 -4724 27852 -4696
rect 27916 -4724 27972 -4696
rect 28036 -4724 28092 -4696
rect 28156 -4724 28212 -4696
rect 28276 -4724 28332 -4696
rect 28396 -4724 28452 -4696
rect 28516 -4724 28572 -4696
rect 28636 -4724 28692 -4696
rect 28756 -4724 28812 -4696
rect 28876 -4724 28932 -4696
rect 28996 -4724 29052 -4696
rect 29116 -4724 29172 -4696
rect 29236 -4724 29292 -4696
rect 29356 -4724 29412 -4696
rect 29476 -4724 29532 -4696
rect 29596 -4724 29652 -4696
rect 29716 -4724 29772 -4696
rect 29836 -4724 29892 -4696
rect 29956 -4724 30012 -4696
rect 30076 -4724 30132 -4696
rect 30196 -4724 30252 -4696
rect 30316 -4724 30372 -4696
rect 30436 -4724 30492 -4696
rect 30556 -4724 30612 -4696
rect 30676 -4724 30732 -4696
rect 30796 -4724 30852 -4696
rect 30916 -4724 30972 -4696
rect 31036 -4724 31092 -4696
rect 31156 -4724 31212 -4696
rect 31276 -4724 31332 -4696
rect 31396 -4724 31452 -4696
rect 31516 -4724 31572 -4696
rect 31636 -4724 31692 -4696
rect 31756 -4724 31812 -4696
rect 31876 -4724 31932 -4696
rect 31996 -4724 32052 -4696
rect 32116 -4724 32172 -4696
rect 32236 -4724 32292 -4696
rect 32356 -4724 32412 -4696
rect 32476 -4724 32532 -4696
rect 32596 -4724 32652 -4696
rect 32716 -4724 32772 -4696
rect 32836 -4724 32892 -4696
rect 32956 -4724 33012 -4696
rect 33076 -4724 33132 -4696
rect 33196 -4724 33252 -4696
rect 33316 -4724 33372 -4696
rect 33436 -4724 33492 -4696
rect 33556 -4724 33612 -4696
rect 33676 -4724 33732 -4696
rect 33796 -4724 33852 -4696
rect 33916 -4724 33972 -4696
rect 34036 -4724 34092 -4696
rect 34156 -4724 34212 -4696
rect 34276 -4724 34332 -4696
rect 34396 -4724 34452 -4696
rect 34516 -4724 34572 -4696
rect 34636 -4724 34692 -4696
rect 34756 -4724 34812 -4696
rect 34876 -4724 34932 -4696
rect 34996 -4724 35052 -4696
rect 35116 -4724 35172 -4696
rect 35236 -4724 35292 -4696
rect 35356 -4724 35412 -4696
rect 35476 -4724 35532 -4696
rect 35596 -4724 35652 -4696
rect 35716 -4724 35772 -4696
rect 35836 -4724 35892 -4696
rect 35956 -4724 36012 -4696
rect 36076 -4724 36132 -4696
rect 36196 -4724 36252 -4696
rect 36316 -4724 36372 -4696
rect 36436 -4724 36492 -4696
rect 36556 -4724 36612 -4696
rect 36676 -4724 36732 -4696
rect 36796 -4724 36852 -4696
rect 36916 -4724 36972 -4696
rect 37036 -4724 37092 -4696
rect 37156 -4724 37212 -4696
rect 37276 -4724 37332 -4696
rect 37396 -4724 37452 -4696
rect 37516 -4724 37572 -4696
rect 37636 -4724 37692 -4696
rect 37756 -4724 37812 -4696
rect 37876 -4724 37932 -4696
rect 37996 -4724 38052 -4696
rect 38116 -4724 38172 -4696
rect 38236 -4724 38292 -4696
rect 38356 -4724 38412 -4696
rect 38476 -4724 38532 -4696
rect 38596 -4724 38652 -4696
rect 38716 -4724 38772 -4696
rect 38836 -4724 38892 -4696
rect 38956 -4724 39012 -4696
rect 39076 -4724 39132 -4696
rect 39196 -4724 39252 -4696
rect 39316 -4724 39372 -4696
rect 39436 -4724 39492 -4696
rect 39556 -4724 39612 -4696
rect 39676 -4724 39732 -4696
rect 39796 -4724 39852 -4696
rect 39916 -4724 39972 -4696
rect 40036 -4724 40092 -4696
rect 40156 -4724 40212 -4696
rect 40276 -4724 40332 -4696
rect 40396 -4724 40452 -4696
rect 40516 -4724 40572 -4696
rect 40636 -4724 40692 -4696
rect 40756 -4724 40812 -4696
rect 40876 -4724 40932 -4696
rect 40996 -4724 41052 -4696
rect 41116 -4724 41172 -4696
rect 41236 -4724 41292 -4696
rect 41356 -4724 41412 -4696
rect 41476 -4724 41532 -4696
rect 41596 -4724 41652 -4696
rect 41716 -4724 41772 -4696
rect 41836 -4724 41892 -4696
rect 41956 -4724 42012 -4696
rect 42076 -4724 42132 -4696
rect 42196 -4724 42252 -4696
rect 42316 -4724 42372 -4696
rect 42436 -4724 42492 -4696
rect 42556 -4724 42612 -4696
rect 42676 -4724 42732 -4696
rect 42796 -4724 42852 -4696
rect 42916 -4724 42972 -4696
rect 43036 -4724 43092 -4696
rect 43156 -4724 43212 -4696
rect 43276 -4724 43332 -4696
rect 43396 -4724 43452 -4696
rect 43516 -4724 43572 -4696
rect 43636 -4724 43692 -4696
rect 43756 -4724 43812 -4696
rect 43876 -4724 43932 -4696
rect 43996 -4724 44052 -4696
rect 44116 -4724 44172 -4696
rect 44236 -4724 44292 -4696
rect 44356 -4724 44412 -4696
rect 44476 -4724 44532 -4696
rect 44596 -4724 44652 -4696
rect 44716 -4724 44772 -4696
rect 44836 -4724 44892 -4696
rect 44956 -4724 45012 -4696
rect 45076 -4724 45132 -4696
rect 45196 -4724 45252 -4696
rect 45316 -4724 45372 -4696
rect 45436 -4724 45492 -4696
rect 45556 -4724 45612 -4696
rect 25848 -4868 25932 -4848
rect 25848 -4876 25868 -4868
rect 25876 -4876 25904 -4868
rect 25912 -4876 25932 -4868
rect 25968 -4868 26052 -4848
rect 25968 -4876 25988 -4868
rect 25996 -4876 26024 -4868
rect 26032 -4876 26052 -4868
rect 26088 -4868 26172 -4848
rect 26088 -4876 26108 -4868
rect 26116 -4876 26144 -4868
rect 26152 -4876 26172 -4868
rect 26208 -4868 26292 -4848
rect 26208 -4876 26228 -4868
rect 26236 -4876 26264 -4868
rect 26272 -4876 26292 -4868
rect 26328 -4868 26412 -4848
rect 26328 -4876 26348 -4868
rect 26356 -4876 26384 -4868
rect 26392 -4876 26412 -4868
rect 26448 -4868 26532 -4848
rect 26448 -4876 26468 -4868
rect 26476 -4876 26504 -4868
rect 26512 -4876 26532 -4868
rect 26568 -4868 26652 -4848
rect 26568 -4876 26588 -4868
rect 26596 -4876 26624 -4868
rect 26632 -4876 26652 -4868
rect 26688 -4868 26772 -4848
rect 26688 -4876 26708 -4868
rect 26716 -4876 26744 -4868
rect 26752 -4876 26772 -4868
rect 26808 -4868 26892 -4848
rect 26808 -4876 26828 -4868
rect 26836 -4876 26864 -4868
rect 26872 -4876 26892 -4868
rect 26928 -4868 27012 -4848
rect 26928 -4876 26948 -4868
rect 26956 -4876 26984 -4868
rect 26992 -4876 27012 -4868
rect 27048 -4868 27132 -4848
rect 27048 -4876 27068 -4868
rect 27076 -4876 27104 -4868
rect 27112 -4876 27132 -4868
rect 27168 -4868 27252 -4848
rect 27168 -4876 27188 -4868
rect 27196 -4876 27224 -4868
rect 27232 -4876 27252 -4868
rect 27288 -4868 27372 -4848
rect 27288 -4876 27308 -4868
rect 27316 -4876 27344 -4868
rect 27352 -4876 27372 -4868
rect 27408 -4868 27492 -4848
rect 27408 -4876 27428 -4868
rect 27436 -4876 27464 -4868
rect 27472 -4876 27492 -4868
rect 27528 -4868 27612 -4848
rect 27528 -4876 27548 -4868
rect 27556 -4876 27584 -4868
rect 27592 -4876 27612 -4868
rect 27648 -4868 27732 -4848
rect 27648 -4876 27668 -4868
rect 27676 -4876 27704 -4868
rect 27712 -4876 27732 -4868
rect 27768 -4868 27852 -4848
rect 27768 -4876 27788 -4868
rect 27796 -4876 27824 -4868
rect 27832 -4876 27852 -4868
rect 27888 -4868 27972 -4848
rect 27888 -4876 27908 -4868
rect 27916 -4876 27944 -4868
rect 27952 -4876 27972 -4868
rect 28008 -4868 28092 -4848
rect 28008 -4876 28028 -4868
rect 28036 -4876 28064 -4868
rect 28072 -4876 28092 -4868
rect 28128 -4868 28212 -4848
rect 28128 -4876 28148 -4868
rect 28156 -4876 28184 -4868
rect 28192 -4876 28212 -4868
rect 28248 -4868 28332 -4848
rect 28248 -4876 28268 -4868
rect 28276 -4876 28304 -4868
rect 28312 -4876 28332 -4868
rect 28368 -4868 28452 -4848
rect 28368 -4876 28388 -4868
rect 28396 -4876 28424 -4868
rect 28432 -4876 28452 -4868
rect 28488 -4868 28572 -4848
rect 28488 -4876 28508 -4868
rect 28516 -4876 28544 -4868
rect 28552 -4876 28572 -4868
rect 28608 -4868 28692 -4848
rect 28608 -4876 28628 -4868
rect 28636 -4876 28664 -4868
rect 28672 -4876 28692 -4868
rect 28728 -4868 28812 -4848
rect 28728 -4876 28748 -4868
rect 28756 -4876 28784 -4868
rect 28792 -4876 28812 -4868
rect 28848 -4868 28932 -4848
rect 28848 -4876 28868 -4868
rect 28876 -4876 28904 -4868
rect 28912 -4876 28932 -4868
rect 28968 -4868 29052 -4848
rect 28968 -4876 28988 -4868
rect 28996 -4876 29024 -4868
rect 29032 -4876 29052 -4868
rect 29088 -4868 29172 -4848
rect 29088 -4876 29108 -4868
rect 29116 -4876 29144 -4868
rect 29152 -4876 29172 -4868
rect 29208 -4868 29292 -4848
rect 29208 -4876 29228 -4868
rect 29236 -4876 29264 -4868
rect 29272 -4876 29292 -4868
rect 29328 -4868 29412 -4848
rect 29328 -4876 29348 -4868
rect 29356 -4876 29384 -4868
rect 29392 -4876 29412 -4868
rect 29448 -4868 29532 -4848
rect 29448 -4876 29468 -4868
rect 29476 -4876 29504 -4868
rect 29512 -4876 29532 -4868
rect 29568 -4868 29652 -4848
rect 29568 -4876 29588 -4868
rect 29596 -4876 29624 -4868
rect 29632 -4876 29652 -4868
rect 29688 -4868 29772 -4848
rect 29688 -4876 29708 -4868
rect 29716 -4876 29744 -4868
rect 29752 -4876 29772 -4868
rect 29808 -4868 29892 -4848
rect 29808 -4876 29828 -4868
rect 29836 -4876 29864 -4868
rect 29872 -4876 29892 -4868
rect 29928 -4868 30012 -4848
rect 29928 -4876 29948 -4868
rect 29956 -4876 29984 -4868
rect 29992 -4876 30012 -4868
rect 30048 -4868 30132 -4848
rect 30048 -4876 30068 -4868
rect 30076 -4876 30104 -4868
rect 30112 -4876 30132 -4868
rect 30168 -4868 30252 -4848
rect 30168 -4876 30188 -4868
rect 30196 -4876 30224 -4868
rect 30232 -4876 30252 -4868
rect 30288 -4868 30372 -4848
rect 30288 -4876 30308 -4868
rect 30316 -4876 30344 -4868
rect 30352 -4876 30372 -4868
rect 30408 -4868 30492 -4848
rect 30408 -4876 30428 -4868
rect 30436 -4876 30464 -4868
rect 30472 -4876 30492 -4868
rect 30528 -4868 30612 -4848
rect 30528 -4876 30548 -4868
rect 30556 -4876 30584 -4868
rect 30592 -4876 30612 -4868
rect 30648 -4868 30732 -4848
rect 30648 -4876 30668 -4868
rect 30676 -4876 30704 -4868
rect 30712 -4876 30732 -4868
rect 30768 -4868 30852 -4848
rect 30768 -4876 30788 -4868
rect 30796 -4876 30824 -4868
rect 30832 -4876 30852 -4868
rect 30888 -4868 30972 -4848
rect 30888 -4876 30908 -4868
rect 30916 -4876 30944 -4868
rect 30952 -4876 30972 -4868
rect 31008 -4868 31092 -4848
rect 31008 -4876 31028 -4868
rect 31036 -4876 31064 -4868
rect 31072 -4876 31092 -4868
rect 31128 -4868 31212 -4848
rect 31128 -4876 31148 -4868
rect 31156 -4876 31184 -4868
rect 31192 -4876 31212 -4868
rect 31248 -4868 31332 -4848
rect 31248 -4876 31268 -4868
rect 31276 -4876 31304 -4868
rect 31312 -4876 31332 -4868
rect 31368 -4868 31452 -4848
rect 31368 -4876 31388 -4868
rect 31396 -4876 31424 -4868
rect 31432 -4876 31452 -4868
rect 31488 -4868 31572 -4848
rect 31488 -4876 31508 -4868
rect 31516 -4876 31544 -4868
rect 31552 -4876 31572 -4868
rect 31608 -4868 31692 -4848
rect 31608 -4876 31628 -4868
rect 31636 -4876 31664 -4868
rect 31672 -4876 31692 -4868
rect 31728 -4868 31812 -4848
rect 31728 -4876 31748 -4868
rect 31756 -4876 31784 -4868
rect 31792 -4876 31812 -4868
rect 31848 -4868 31932 -4848
rect 31848 -4876 31868 -4868
rect 31876 -4876 31904 -4868
rect 31912 -4876 31932 -4868
rect 31968 -4868 32052 -4848
rect 31968 -4876 31988 -4868
rect 31996 -4876 32024 -4868
rect 32032 -4876 32052 -4868
rect 32088 -4868 32172 -4848
rect 32088 -4876 32108 -4868
rect 32116 -4876 32144 -4868
rect 32152 -4876 32172 -4868
rect 32208 -4868 32292 -4848
rect 32208 -4876 32228 -4868
rect 32236 -4876 32264 -4868
rect 32272 -4876 32292 -4868
rect 32328 -4868 32412 -4848
rect 32328 -4876 32348 -4868
rect 32356 -4876 32384 -4868
rect 32392 -4876 32412 -4868
rect 32448 -4868 32532 -4848
rect 32448 -4876 32468 -4868
rect 32476 -4876 32504 -4868
rect 32512 -4876 32532 -4868
rect 32568 -4868 32652 -4848
rect 32568 -4876 32588 -4868
rect 32596 -4876 32624 -4868
rect 32632 -4876 32652 -4868
rect 32688 -4868 32772 -4848
rect 32688 -4876 32708 -4868
rect 32716 -4876 32744 -4868
rect 32752 -4876 32772 -4868
rect 32808 -4868 32892 -4848
rect 32808 -4876 32828 -4868
rect 32836 -4876 32864 -4868
rect 32872 -4876 32892 -4868
rect 32928 -4868 33012 -4848
rect 32928 -4876 32948 -4868
rect 32956 -4876 32984 -4868
rect 32992 -4876 33012 -4868
rect 33048 -4868 33132 -4848
rect 33048 -4876 33068 -4868
rect 33076 -4876 33104 -4868
rect 33112 -4876 33132 -4868
rect 33168 -4868 33252 -4848
rect 33168 -4876 33188 -4868
rect 33196 -4876 33224 -4868
rect 33232 -4876 33252 -4868
rect 33288 -4868 33372 -4848
rect 33288 -4876 33308 -4868
rect 33316 -4876 33344 -4868
rect 33352 -4876 33372 -4868
rect 33408 -4868 33492 -4848
rect 33408 -4876 33428 -4868
rect 33436 -4876 33464 -4868
rect 33472 -4876 33492 -4868
rect 33528 -4868 33612 -4848
rect 33528 -4876 33548 -4868
rect 33556 -4876 33584 -4868
rect 33592 -4876 33612 -4868
rect 33648 -4868 33732 -4848
rect 33648 -4876 33668 -4868
rect 33676 -4876 33704 -4868
rect 33712 -4876 33732 -4868
rect 33768 -4868 33852 -4848
rect 33768 -4876 33788 -4868
rect 33796 -4876 33824 -4868
rect 33832 -4876 33852 -4868
rect 33888 -4868 33972 -4848
rect 33888 -4876 33908 -4868
rect 33916 -4876 33944 -4868
rect 33952 -4876 33972 -4868
rect 34008 -4868 34092 -4848
rect 34008 -4876 34028 -4868
rect 34036 -4876 34064 -4868
rect 34072 -4876 34092 -4868
rect 34128 -4868 34212 -4848
rect 34128 -4876 34148 -4868
rect 34156 -4876 34184 -4868
rect 34192 -4876 34212 -4868
rect 34248 -4868 34332 -4848
rect 34248 -4876 34268 -4868
rect 34276 -4876 34304 -4868
rect 34312 -4876 34332 -4868
rect 34368 -4868 34452 -4848
rect 34368 -4876 34388 -4868
rect 34396 -4876 34424 -4868
rect 34432 -4876 34452 -4868
rect 34488 -4868 34572 -4848
rect 34488 -4876 34508 -4868
rect 34516 -4876 34544 -4868
rect 34552 -4876 34572 -4868
rect 34608 -4868 34692 -4848
rect 34608 -4876 34628 -4868
rect 34636 -4876 34664 -4868
rect 34672 -4876 34692 -4868
rect 34728 -4868 34812 -4848
rect 34728 -4876 34748 -4868
rect 34756 -4876 34784 -4868
rect 34792 -4876 34812 -4868
rect 34848 -4868 34932 -4848
rect 34848 -4876 34868 -4868
rect 34876 -4876 34904 -4868
rect 34912 -4876 34932 -4868
rect 34968 -4868 35052 -4848
rect 34968 -4876 34988 -4868
rect 34996 -4876 35024 -4868
rect 35032 -4876 35052 -4868
rect 35088 -4868 35172 -4848
rect 35088 -4876 35108 -4868
rect 35116 -4876 35144 -4868
rect 35152 -4876 35172 -4868
rect 35208 -4868 35292 -4848
rect 35208 -4876 35228 -4868
rect 35236 -4876 35264 -4868
rect 35272 -4876 35292 -4868
rect 35328 -4868 35412 -4848
rect 35328 -4876 35348 -4868
rect 35356 -4876 35384 -4868
rect 35392 -4876 35412 -4868
rect 35448 -4868 35532 -4848
rect 35448 -4876 35468 -4868
rect 35476 -4876 35504 -4868
rect 35512 -4876 35532 -4868
rect 35568 -4868 35652 -4848
rect 35568 -4876 35588 -4868
rect 35596 -4876 35624 -4868
rect 35632 -4876 35652 -4868
rect 35688 -4868 35772 -4848
rect 35688 -4876 35708 -4868
rect 35716 -4876 35744 -4868
rect 35752 -4876 35772 -4868
rect 35808 -4868 35892 -4848
rect 35808 -4876 35828 -4868
rect 35836 -4876 35864 -4868
rect 35872 -4876 35892 -4868
rect 35928 -4868 36012 -4848
rect 35928 -4876 35948 -4868
rect 35956 -4876 35984 -4868
rect 35992 -4876 36012 -4868
rect 36048 -4868 36132 -4848
rect 36048 -4876 36068 -4868
rect 36076 -4876 36104 -4868
rect 36112 -4876 36132 -4868
rect 36168 -4868 36252 -4848
rect 36168 -4876 36188 -4868
rect 36196 -4876 36224 -4868
rect 36232 -4876 36252 -4868
rect 36288 -4868 36372 -4848
rect 36288 -4876 36308 -4868
rect 36316 -4876 36344 -4868
rect 36352 -4876 36372 -4868
rect 36408 -4868 36492 -4848
rect 36408 -4876 36428 -4868
rect 36436 -4876 36464 -4868
rect 36472 -4876 36492 -4868
rect 36528 -4868 36612 -4848
rect 36528 -4876 36548 -4868
rect 36556 -4876 36584 -4868
rect 36592 -4876 36612 -4868
rect 36648 -4868 36732 -4848
rect 36648 -4876 36668 -4868
rect 36676 -4876 36704 -4868
rect 36712 -4876 36732 -4868
rect 36768 -4868 36852 -4848
rect 36768 -4876 36788 -4868
rect 36796 -4876 36824 -4868
rect 36832 -4876 36852 -4868
rect 36888 -4868 36972 -4848
rect 36888 -4876 36908 -4868
rect 36916 -4876 36944 -4868
rect 36952 -4876 36972 -4868
rect 37008 -4868 37092 -4848
rect 37008 -4876 37028 -4868
rect 37036 -4876 37064 -4868
rect 37072 -4876 37092 -4868
rect 37128 -4868 37212 -4848
rect 37128 -4876 37148 -4868
rect 37156 -4876 37184 -4868
rect 37192 -4876 37212 -4868
rect 37248 -4868 37332 -4848
rect 37248 -4876 37268 -4868
rect 37276 -4876 37304 -4868
rect 37312 -4876 37332 -4868
rect 37368 -4868 37452 -4848
rect 37368 -4876 37388 -4868
rect 37396 -4876 37424 -4868
rect 37432 -4876 37452 -4868
rect 37488 -4868 37572 -4848
rect 37488 -4876 37508 -4868
rect 37516 -4876 37544 -4868
rect 37552 -4876 37572 -4868
rect 37608 -4868 37692 -4848
rect 37608 -4876 37628 -4868
rect 37636 -4876 37664 -4868
rect 37672 -4876 37692 -4868
rect 37728 -4868 37812 -4848
rect 37728 -4876 37748 -4868
rect 37756 -4876 37784 -4868
rect 37792 -4876 37812 -4868
rect 37848 -4868 37932 -4848
rect 37848 -4876 37868 -4868
rect 37876 -4876 37904 -4868
rect 37912 -4876 37932 -4868
rect 37968 -4868 38052 -4848
rect 37968 -4876 37988 -4868
rect 37996 -4876 38024 -4868
rect 38032 -4876 38052 -4868
rect 38088 -4868 38172 -4848
rect 38088 -4876 38108 -4868
rect 38116 -4876 38144 -4868
rect 38152 -4876 38172 -4868
rect 38208 -4868 38292 -4848
rect 38208 -4876 38228 -4868
rect 38236 -4876 38264 -4868
rect 38272 -4876 38292 -4868
rect 38328 -4868 38412 -4848
rect 38328 -4876 38348 -4868
rect 38356 -4876 38384 -4868
rect 38392 -4876 38412 -4868
rect 38448 -4868 38532 -4848
rect 38448 -4876 38468 -4868
rect 38476 -4876 38504 -4868
rect 38512 -4876 38532 -4868
rect 38568 -4868 38652 -4848
rect 38568 -4876 38588 -4868
rect 38596 -4876 38624 -4868
rect 38632 -4876 38652 -4868
rect 38688 -4868 38772 -4848
rect 38688 -4876 38708 -4868
rect 38716 -4876 38744 -4868
rect 38752 -4876 38772 -4868
rect 38808 -4868 38892 -4848
rect 38808 -4876 38828 -4868
rect 38836 -4876 38864 -4868
rect 38872 -4876 38892 -4868
rect 38928 -4868 39012 -4848
rect 38928 -4876 38948 -4868
rect 38956 -4876 38984 -4868
rect 38992 -4876 39012 -4868
rect 39048 -4868 39132 -4848
rect 39048 -4876 39068 -4868
rect 39076 -4876 39104 -4868
rect 39112 -4876 39132 -4868
rect 39168 -4868 39252 -4848
rect 39168 -4876 39188 -4868
rect 39196 -4876 39224 -4868
rect 39232 -4876 39252 -4868
rect 39288 -4868 39372 -4848
rect 39288 -4876 39308 -4868
rect 39316 -4876 39344 -4868
rect 39352 -4876 39372 -4868
rect 39408 -4868 39492 -4848
rect 39408 -4876 39428 -4868
rect 39436 -4876 39464 -4868
rect 39472 -4876 39492 -4868
rect 39528 -4868 39612 -4848
rect 39528 -4876 39548 -4868
rect 39556 -4876 39584 -4868
rect 39592 -4876 39612 -4868
rect 39648 -4868 39732 -4848
rect 39648 -4876 39668 -4868
rect 39676 -4876 39704 -4868
rect 39712 -4876 39732 -4868
rect 39768 -4868 39852 -4848
rect 39768 -4876 39788 -4868
rect 39796 -4876 39824 -4868
rect 39832 -4876 39852 -4868
rect 39888 -4868 39972 -4848
rect 39888 -4876 39908 -4868
rect 39916 -4876 39944 -4868
rect 39952 -4876 39972 -4868
rect 40008 -4868 40092 -4848
rect 40008 -4876 40028 -4868
rect 40036 -4876 40064 -4868
rect 40072 -4876 40092 -4868
rect 40128 -4868 40212 -4848
rect 40128 -4876 40148 -4868
rect 40156 -4876 40184 -4868
rect 40192 -4876 40212 -4868
rect 40248 -4868 40332 -4848
rect 40248 -4876 40268 -4868
rect 40276 -4876 40304 -4868
rect 40312 -4876 40332 -4868
rect 40368 -4868 40452 -4848
rect 40368 -4876 40388 -4868
rect 40396 -4876 40424 -4868
rect 40432 -4876 40452 -4868
rect 40488 -4868 40572 -4848
rect 40488 -4876 40508 -4868
rect 40516 -4876 40544 -4868
rect 40552 -4876 40572 -4868
rect 40608 -4868 40692 -4848
rect 40608 -4876 40628 -4868
rect 40636 -4876 40664 -4868
rect 40672 -4876 40692 -4868
rect 40728 -4868 40812 -4848
rect 40728 -4876 40748 -4868
rect 40756 -4876 40784 -4868
rect 40792 -4876 40812 -4868
rect 40848 -4868 40932 -4848
rect 40848 -4876 40868 -4868
rect 40876 -4876 40904 -4868
rect 40912 -4876 40932 -4868
rect 40968 -4868 41052 -4848
rect 40968 -4876 40988 -4868
rect 40996 -4876 41024 -4868
rect 41032 -4876 41052 -4868
rect 41088 -4868 41172 -4848
rect 41088 -4876 41108 -4868
rect 41116 -4876 41144 -4868
rect 41152 -4876 41172 -4868
rect 41208 -4868 41292 -4848
rect 41208 -4876 41228 -4868
rect 41236 -4876 41264 -4868
rect 41272 -4876 41292 -4868
rect 41328 -4868 41412 -4848
rect 41328 -4876 41348 -4868
rect 41356 -4876 41384 -4868
rect 41392 -4876 41412 -4868
rect 41448 -4868 41532 -4848
rect 41448 -4876 41468 -4868
rect 41476 -4876 41504 -4868
rect 41512 -4876 41532 -4868
rect 41568 -4868 41652 -4848
rect 41568 -4876 41588 -4868
rect 41596 -4876 41624 -4868
rect 41632 -4876 41652 -4868
rect 41688 -4868 41772 -4848
rect 41688 -4876 41708 -4868
rect 41716 -4876 41744 -4868
rect 41752 -4876 41772 -4868
rect 41808 -4868 41892 -4848
rect 41808 -4876 41828 -4868
rect 41836 -4876 41864 -4868
rect 41872 -4876 41892 -4868
rect 41928 -4868 42012 -4848
rect 41928 -4876 41948 -4868
rect 41956 -4876 41984 -4868
rect 41992 -4876 42012 -4868
rect 42048 -4868 42132 -4848
rect 42048 -4876 42068 -4868
rect 42076 -4876 42104 -4868
rect 42112 -4876 42132 -4868
rect 42168 -4868 42252 -4848
rect 42168 -4876 42188 -4868
rect 42196 -4876 42224 -4868
rect 42232 -4876 42252 -4868
rect 42288 -4868 42372 -4848
rect 42288 -4876 42308 -4868
rect 42316 -4876 42344 -4868
rect 42352 -4876 42372 -4868
rect 42408 -4868 42492 -4848
rect 42408 -4876 42428 -4868
rect 42436 -4876 42464 -4868
rect 42472 -4876 42492 -4868
rect 42528 -4868 42612 -4848
rect 42528 -4876 42548 -4868
rect 42556 -4876 42584 -4868
rect 42592 -4876 42612 -4868
rect 42648 -4868 42732 -4848
rect 42648 -4876 42668 -4868
rect 42676 -4876 42704 -4868
rect 42712 -4876 42732 -4868
rect 42768 -4868 42852 -4848
rect 42768 -4876 42788 -4868
rect 42796 -4876 42824 -4868
rect 42832 -4876 42852 -4868
rect 42888 -4868 42972 -4848
rect 42888 -4876 42908 -4868
rect 42916 -4876 42944 -4868
rect 42952 -4876 42972 -4868
rect 43008 -4868 43092 -4848
rect 43008 -4876 43028 -4868
rect 43036 -4876 43064 -4868
rect 43072 -4876 43092 -4868
rect 43128 -4868 43212 -4848
rect 43128 -4876 43148 -4868
rect 43156 -4876 43184 -4868
rect 43192 -4876 43212 -4868
rect 43248 -4868 43332 -4848
rect 43248 -4876 43268 -4868
rect 43276 -4876 43304 -4868
rect 43312 -4876 43332 -4868
rect 43368 -4868 43452 -4848
rect 43368 -4876 43388 -4868
rect 43396 -4876 43424 -4868
rect 43432 -4876 43452 -4868
rect 43488 -4868 43572 -4848
rect 43488 -4876 43508 -4868
rect 43516 -4876 43544 -4868
rect 43552 -4876 43572 -4868
rect 43608 -4868 43692 -4848
rect 43608 -4876 43628 -4868
rect 43636 -4876 43664 -4868
rect 43672 -4876 43692 -4868
rect 43728 -4868 43812 -4848
rect 43728 -4876 43748 -4868
rect 43756 -4876 43784 -4868
rect 43792 -4876 43812 -4868
rect 43848 -4868 43932 -4848
rect 43848 -4876 43868 -4868
rect 43876 -4876 43904 -4868
rect 43912 -4876 43932 -4868
rect 43968 -4868 44052 -4848
rect 43968 -4876 43988 -4868
rect 43996 -4876 44024 -4868
rect 44032 -4876 44052 -4868
rect 44088 -4868 44172 -4848
rect 44088 -4876 44108 -4868
rect 44116 -4876 44144 -4868
rect 44152 -4876 44172 -4868
rect 44208 -4868 44292 -4848
rect 44208 -4876 44228 -4868
rect 44236 -4876 44264 -4868
rect 44272 -4876 44292 -4868
rect 44328 -4868 44412 -4848
rect 44328 -4876 44348 -4868
rect 44356 -4876 44384 -4868
rect 44392 -4876 44412 -4868
rect 44448 -4868 44532 -4848
rect 44448 -4876 44468 -4868
rect 44476 -4876 44504 -4868
rect 44512 -4876 44532 -4868
rect 44568 -4868 44652 -4848
rect 44568 -4876 44588 -4868
rect 44596 -4876 44624 -4868
rect 44632 -4876 44652 -4868
rect 44688 -4868 44772 -4848
rect 44688 -4876 44708 -4868
rect 44716 -4876 44744 -4868
rect 44752 -4876 44772 -4868
rect 44808 -4868 44892 -4848
rect 44808 -4876 44828 -4868
rect 44836 -4876 44864 -4868
rect 44872 -4876 44892 -4868
rect 44928 -4868 45012 -4848
rect 44928 -4876 44948 -4868
rect 44956 -4876 44984 -4868
rect 44992 -4876 45012 -4868
rect 45048 -4868 45132 -4848
rect 45048 -4876 45068 -4868
rect 45076 -4876 45104 -4868
rect 45112 -4876 45132 -4868
rect 45168 -4868 45252 -4848
rect 45168 -4876 45188 -4868
rect 45196 -4876 45224 -4868
rect 45232 -4876 45252 -4868
rect 45288 -4868 45372 -4848
rect 45288 -4876 45308 -4868
rect 45316 -4876 45344 -4868
rect 45352 -4876 45372 -4868
rect 45408 -4868 45492 -4848
rect 45408 -4876 45428 -4868
rect 45436 -4876 45464 -4868
rect 45472 -4876 45492 -4868
rect 45528 -4868 45612 -4848
rect 45528 -4876 45548 -4868
rect 45556 -4876 45584 -4868
rect 45592 -4876 45612 -4868
rect 25876 -4904 25932 -4876
rect 25996 -4904 26052 -4876
rect 26116 -4904 26172 -4876
rect 26236 -4904 26292 -4876
rect 26356 -4904 26412 -4876
rect 26476 -4904 26532 -4876
rect 26596 -4904 26652 -4876
rect 26716 -4904 26772 -4876
rect 26836 -4904 26892 -4876
rect 26956 -4904 27012 -4876
rect 27076 -4904 27132 -4876
rect 27196 -4904 27252 -4876
rect 27316 -4904 27372 -4876
rect 27436 -4904 27492 -4876
rect 27556 -4904 27612 -4876
rect 27676 -4904 27732 -4876
rect 27796 -4904 27852 -4876
rect 27916 -4904 27972 -4876
rect 28036 -4904 28092 -4876
rect 28156 -4904 28212 -4876
rect 28276 -4904 28332 -4876
rect 28396 -4904 28452 -4876
rect 28516 -4904 28572 -4876
rect 28636 -4904 28692 -4876
rect 28756 -4904 28812 -4876
rect 28876 -4904 28932 -4876
rect 28996 -4904 29052 -4876
rect 29116 -4904 29172 -4876
rect 29236 -4904 29292 -4876
rect 29356 -4904 29412 -4876
rect 29476 -4904 29532 -4876
rect 29596 -4904 29652 -4876
rect 29716 -4904 29772 -4876
rect 29836 -4904 29892 -4876
rect 29956 -4904 30012 -4876
rect 30076 -4904 30132 -4876
rect 30196 -4904 30252 -4876
rect 30316 -4904 30372 -4876
rect 30436 -4904 30492 -4876
rect 30556 -4904 30612 -4876
rect 30676 -4904 30732 -4876
rect 30796 -4904 30852 -4876
rect 30916 -4904 30972 -4876
rect 31036 -4904 31092 -4876
rect 31156 -4904 31212 -4876
rect 31276 -4904 31332 -4876
rect 31396 -4904 31452 -4876
rect 31516 -4904 31572 -4876
rect 31636 -4904 31692 -4876
rect 31756 -4904 31812 -4876
rect 31876 -4904 31932 -4876
rect 31996 -4904 32052 -4876
rect 32116 -4904 32172 -4876
rect 32236 -4904 32292 -4876
rect 32356 -4904 32412 -4876
rect 32476 -4904 32532 -4876
rect 32596 -4904 32652 -4876
rect 32716 -4904 32772 -4876
rect 32836 -4904 32892 -4876
rect 32956 -4904 33012 -4876
rect 33076 -4904 33132 -4876
rect 33196 -4904 33252 -4876
rect 33316 -4904 33372 -4876
rect 33436 -4904 33492 -4876
rect 33556 -4904 33612 -4876
rect 33676 -4904 33732 -4876
rect 33796 -4904 33852 -4876
rect 33916 -4904 33972 -4876
rect 34036 -4904 34092 -4876
rect 34156 -4904 34212 -4876
rect 34276 -4904 34332 -4876
rect 34396 -4904 34452 -4876
rect 34516 -4904 34572 -4876
rect 34636 -4904 34692 -4876
rect 34756 -4904 34812 -4876
rect 34876 -4904 34932 -4876
rect 34996 -4904 35052 -4876
rect 35116 -4904 35172 -4876
rect 35236 -4904 35292 -4876
rect 35356 -4904 35412 -4876
rect 35476 -4904 35532 -4876
rect 35596 -4904 35652 -4876
rect 35716 -4904 35772 -4876
rect 35836 -4904 35892 -4876
rect 35956 -4904 36012 -4876
rect 36076 -4904 36132 -4876
rect 36196 -4904 36252 -4876
rect 36316 -4904 36372 -4876
rect 36436 -4904 36492 -4876
rect 36556 -4904 36612 -4876
rect 36676 -4904 36732 -4876
rect 36796 -4904 36852 -4876
rect 36916 -4904 36972 -4876
rect 37036 -4904 37092 -4876
rect 37156 -4904 37212 -4876
rect 37276 -4904 37332 -4876
rect 37396 -4904 37452 -4876
rect 37516 -4904 37572 -4876
rect 37636 -4904 37692 -4876
rect 37756 -4904 37812 -4876
rect 37876 -4904 37932 -4876
rect 37996 -4904 38052 -4876
rect 38116 -4904 38172 -4876
rect 38236 -4904 38292 -4876
rect 38356 -4904 38412 -4876
rect 38476 -4904 38532 -4876
rect 38596 -4904 38652 -4876
rect 38716 -4904 38772 -4876
rect 38836 -4904 38892 -4876
rect 38956 -4904 39012 -4876
rect 39076 -4904 39132 -4876
rect 39196 -4904 39252 -4876
rect 39316 -4904 39372 -4876
rect 39436 -4904 39492 -4876
rect 39556 -4904 39612 -4876
rect 39676 -4904 39732 -4876
rect 39796 -4904 39852 -4876
rect 39916 -4904 39972 -4876
rect 40036 -4904 40092 -4876
rect 40156 -4904 40212 -4876
rect 40276 -4904 40332 -4876
rect 40396 -4904 40452 -4876
rect 40516 -4904 40572 -4876
rect 40636 -4904 40692 -4876
rect 40756 -4904 40812 -4876
rect 40876 -4904 40932 -4876
rect 40996 -4904 41052 -4876
rect 41116 -4904 41172 -4876
rect 41236 -4904 41292 -4876
rect 41356 -4904 41412 -4876
rect 41476 -4904 41532 -4876
rect 41596 -4904 41652 -4876
rect 41716 -4904 41772 -4876
rect 41836 -4904 41892 -4876
rect 41956 -4904 42012 -4876
rect 42076 -4904 42132 -4876
rect 42196 -4904 42252 -4876
rect 42316 -4904 42372 -4876
rect 42436 -4904 42492 -4876
rect 42556 -4904 42612 -4876
rect 42676 -4904 42732 -4876
rect 42796 -4904 42852 -4876
rect 42916 -4904 42972 -4876
rect 43036 -4904 43092 -4876
rect 43156 -4904 43212 -4876
rect 43276 -4904 43332 -4876
rect 43396 -4904 43452 -4876
rect 43516 -4904 43572 -4876
rect 43636 -4904 43692 -4876
rect 43756 -4904 43812 -4876
rect 43876 -4904 43932 -4876
rect 43996 -4904 44052 -4876
rect 44116 -4904 44172 -4876
rect 44236 -4904 44292 -4876
rect 44356 -4904 44412 -4876
rect 44476 -4904 44532 -4876
rect 44596 -4904 44652 -4876
rect 44716 -4904 44772 -4876
rect 44836 -4904 44892 -4876
rect 44956 -4904 45012 -4876
rect 45076 -4904 45132 -4876
rect 45196 -4904 45252 -4876
rect 45316 -4904 45372 -4876
rect 45436 -4904 45492 -4876
rect 45556 -4904 45612 -4876
rect 25848 -6368 25932 -6348
rect 25848 -6376 25868 -6368
rect 25876 -6376 25904 -6368
rect 25912 -6376 25932 -6368
rect 26088 -6368 26172 -6348
rect 26088 -6376 26108 -6368
rect 26116 -6376 26144 -6368
rect 26152 -6376 26172 -6368
rect 26208 -6368 26292 -6348
rect 26208 -6376 26228 -6368
rect 26236 -6376 26264 -6368
rect 26272 -6376 26292 -6368
rect 26448 -6368 26532 -6348
rect 26448 -6376 26468 -6368
rect 26476 -6376 26504 -6368
rect 26512 -6376 26532 -6368
rect 26568 -6368 26652 -6348
rect 26568 -6376 26588 -6368
rect 26596 -6376 26624 -6368
rect 26632 -6376 26652 -6368
rect 26808 -6368 26892 -6348
rect 26808 -6376 26828 -6368
rect 26836 -6376 26864 -6368
rect 26872 -6376 26892 -6368
rect 26928 -6368 27012 -6348
rect 26928 -6376 26948 -6368
rect 26956 -6376 26984 -6368
rect 26992 -6376 27012 -6368
rect 27168 -6368 27252 -6348
rect 27168 -6376 27188 -6368
rect 27196 -6376 27224 -6368
rect 27232 -6376 27252 -6368
rect 27288 -6368 27372 -6348
rect 27288 -6376 27308 -6368
rect 27316 -6376 27344 -6368
rect 27352 -6376 27372 -6368
rect 27528 -6368 27612 -6348
rect 27528 -6376 27548 -6368
rect 27556 -6376 27584 -6368
rect 27592 -6376 27612 -6368
rect 27648 -6368 27732 -6348
rect 27648 -6376 27668 -6368
rect 27676 -6376 27704 -6368
rect 27712 -6376 27732 -6368
rect 27888 -6368 27972 -6348
rect 27888 -6376 27908 -6368
rect 27916 -6376 27944 -6368
rect 27952 -6376 27972 -6368
rect 28008 -6368 28092 -6348
rect 28008 -6376 28028 -6368
rect 28036 -6376 28064 -6368
rect 28072 -6376 28092 -6368
rect 28248 -6368 28332 -6348
rect 28248 -6376 28268 -6368
rect 28276 -6376 28304 -6368
rect 28312 -6376 28332 -6368
rect 28368 -6368 28452 -6348
rect 28368 -6376 28388 -6368
rect 28396 -6376 28424 -6368
rect 28432 -6376 28452 -6368
rect 28608 -6368 28692 -6348
rect 28608 -6376 28628 -6368
rect 28636 -6376 28664 -6368
rect 28672 -6376 28692 -6368
rect 28728 -6368 28812 -6348
rect 28728 -6376 28748 -6368
rect 28756 -6376 28784 -6368
rect 28792 -6376 28812 -6368
rect 28968 -6368 29052 -6348
rect 28968 -6376 28988 -6368
rect 28996 -6376 29024 -6368
rect 29032 -6376 29052 -6368
rect 29088 -6368 29172 -6348
rect 29088 -6376 29108 -6368
rect 29116 -6376 29144 -6368
rect 29152 -6376 29172 -6368
rect 29328 -6368 29412 -6348
rect 29328 -6376 29348 -6368
rect 29356 -6376 29384 -6368
rect 29392 -6376 29412 -6368
rect 29448 -6368 29532 -6348
rect 29448 -6376 29468 -6368
rect 29476 -6376 29504 -6368
rect 29512 -6376 29532 -6368
rect 29688 -6368 29772 -6348
rect 29688 -6376 29708 -6368
rect 29716 -6376 29744 -6368
rect 29752 -6376 29772 -6368
rect 29808 -6368 29892 -6348
rect 29808 -6376 29828 -6368
rect 29836 -6376 29864 -6368
rect 29872 -6376 29892 -6368
rect 30048 -6368 30132 -6348
rect 30048 -6376 30068 -6368
rect 30076 -6376 30104 -6368
rect 30112 -6376 30132 -6368
rect 30168 -6368 30252 -6348
rect 30168 -6376 30188 -6368
rect 30196 -6376 30224 -6368
rect 30232 -6376 30252 -6368
rect 30408 -6368 30492 -6348
rect 30408 -6376 30428 -6368
rect 30436 -6376 30464 -6368
rect 30472 -6376 30492 -6368
rect 30528 -6368 30612 -6348
rect 30528 -6376 30548 -6368
rect 30556 -6376 30584 -6368
rect 30592 -6376 30612 -6368
rect 30768 -6368 30852 -6348
rect 30768 -6376 30788 -6368
rect 30796 -6376 30824 -6368
rect 30832 -6376 30852 -6368
rect 30888 -6368 30972 -6348
rect 30888 -6376 30908 -6368
rect 30916 -6376 30944 -6368
rect 30952 -6376 30972 -6368
rect 31128 -6368 31212 -6348
rect 31128 -6376 31148 -6368
rect 31156 -6376 31184 -6368
rect 31192 -6376 31212 -6368
rect 31248 -6368 31332 -6348
rect 31248 -6376 31268 -6368
rect 31276 -6376 31304 -6368
rect 31312 -6376 31332 -6368
rect 31488 -6368 31572 -6348
rect 31488 -6376 31508 -6368
rect 31516 -6376 31544 -6368
rect 31552 -6376 31572 -6368
rect 31608 -6368 31692 -6348
rect 31608 -6376 31628 -6368
rect 31636 -6376 31664 -6368
rect 31672 -6376 31692 -6368
rect 31848 -6368 31932 -6348
rect 31848 -6376 31868 -6368
rect 31876 -6376 31904 -6368
rect 31912 -6376 31932 -6368
rect 31968 -6368 32052 -6348
rect 31968 -6376 31988 -6368
rect 31996 -6376 32024 -6368
rect 32032 -6376 32052 -6368
rect 32208 -6368 32292 -6348
rect 32208 -6376 32228 -6368
rect 32236 -6376 32264 -6368
rect 32272 -6376 32292 -6368
rect 32328 -6368 32412 -6348
rect 32328 -6376 32348 -6368
rect 32356 -6376 32384 -6368
rect 32392 -6376 32412 -6368
rect 32568 -6368 32652 -6348
rect 32568 -6376 32588 -6368
rect 32596 -6376 32624 -6368
rect 32632 -6376 32652 -6368
rect 32688 -6368 32772 -6348
rect 32688 -6376 32708 -6368
rect 32716 -6376 32744 -6368
rect 32752 -6376 32772 -6368
rect 32928 -6368 33012 -6348
rect 32928 -6376 32948 -6368
rect 32956 -6376 32984 -6368
rect 32992 -6376 33012 -6368
rect 33048 -6368 33132 -6348
rect 33048 -6376 33068 -6368
rect 33076 -6376 33104 -6368
rect 33112 -6376 33132 -6368
rect 33288 -6368 33372 -6348
rect 33288 -6376 33308 -6368
rect 33316 -6376 33344 -6368
rect 33352 -6376 33372 -6368
rect 33408 -6368 33492 -6348
rect 33408 -6376 33428 -6368
rect 33436 -6376 33464 -6368
rect 33472 -6376 33492 -6368
rect 33648 -6368 33732 -6348
rect 33648 -6376 33668 -6368
rect 33676 -6376 33704 -6368
rect 33712 -6376 33732 -6368
rect 33768 -6368 33852 -6348
rect 33768 -6376 33788 -6368
rect 33796 -6376 33824 -6368
rect 33832 -6376 33852 -6368
rect 34008 -6368 34092 -6348
rect 34008 -6376 34028 -6368
rect 34036 -6376 34064 -6368
rect 34072 -6376 34092 -6368
rect 34128 -6368 34212 -6348
rect 34128 -6376 34148 -6368
rect 34156 -6376 34184 -6368
rect 34192 -6376 34212 -6368
rect 34368 -6368 34452 -6348
rect 34368 -6376 34388 -6368
rect 34396 -6376 34424 -6368
rect 34432 -6376 34452 -6368
rect 34488 -6368 34572 -6348
rect 34488 -6376 34508 -6368
rect 34516 -6376 34544 -6368
rect 34552 -6376 34572 -6368
rect 34728 -6368 34812 -6348
rect 34728 -6376 34748 -6368
rect 34756 -6376 34784 -6368
rect 34792 -6376 34812 -6368
rect 34848 -6368 34932 -6348
rect 34848 -6376 34868 -6368
rect 34876 -6376 34904 -6368
rect 34912 -6376 34932 -6368
rect 35088 -6368 35172 -6348
rect 35088 -6376 35108 -6368
rect 35116 -6376 35144 -6368
rect 35152 -6376 35172 -6368
rect 35208 -6368 35292 -6348
rect 35208 -6376 35228 -6368
rect 35236 -6376 35264 -6368
rect 35272 -6376 35292 -6368
rect 35448 -6368 35532 -6348
rect 35448 -6376 35468 -6368
rect 35476 -6376 35504 -6368
rect 35512 -6376 35532 -6368
rect 35568 -6368 35652 -6348
rect 35568 -6376 35588 -6368
rect 35596 -6376 35624 -6368
rect 35632 -6376 35652 -6368
rect 35808 -6368 35892 -6348
rect 35808 -6376 35828 -6368
rect 35836 -6376 35864 -6368
rect 35872 -6376 35892 -6368
rect 35928 -6368 36012 -6348
rect 35928 -6376 35948 -6368
rect 35956 -6376 35984 -6368
rect 35992 -6376 36012 -6368
rect 36168 -6368 36252 -6348
rect 36168 -6376 36188 -6368
rect 36196 -6376 36224 -6368
rect 36232 -6376 36252 -6368
rect 36288 -6368 36372 -6348
rect 36288 -6376 36308 -6368
rect 36316 -6376 36344 -6368
rect 36352 -6376 36372 -6368
rect 36528 -6368 36612 -6348
rect 36528 -6376 36548 -6368
rect 36556 -6376 36584 -6368
rect 36592 -6376 36612 -6368
rect 36648 -6368 36732 -6348
rect 36648 -6376 36668 -6368
rect 36676 -6376 36704 -6368
rect 36712 -6376 36732 -6368
rect 36888 -6368 36972 -6348
rect 36888 -6376 36908 -6368
rect 36916 -6376 36944 -6368
rect 36952 -6376 36972 -6368
rect 37008 -6368 37092 -6348
rect 37008 -6376 37028 -6368
rect 37036 -6376 37064 -6368
rect 37072 -6376 37092 -6368
rect 37248 -6368 37332 -6348
rect 37248 -6376 37268 -6368
rect 37276 -6376 37304 -6368
rect 37312 -6376 37332 -6368
rect 37368 -6368 37452 -6348
rect 37368 -6376 37388 -6368
rect 37396 -6376 37424 -6368
rect 37432 -6376 37452 -6368
rect 37608 -6368 37692 -6348
rect 37608 -6376 37628 -6368
rect 37636 -6376 37664 -6368
rect 37672 -6376 37692 -6368
rect 37728 -6368 37812 -6348
rect 37728 -6376 37748 -6368
rect 37756 -6376 37784 -6368
rect 37792 -6376 37812 -6368
rect 37968 -6368 38052 -6348
rect 37968 -6376 37988 -6368
rect 37996 -6376 38024 -6368
rect 38032 -6376 38052 -6368
rect 38088 -6368 38172 -6348
rect 38088 -6376 38108 -6368
rect 38116 -6376 38144 -6368
rect 38152 -6376 38172 -6368
rect 38328 -6368 38412 -6348
rect 38328 -6376 38348 -6368
rect 38356 -6376 38384 -6368
rect 38392 -6376 38412 -6368
rect 38448 -6368 38532 -6348
rect 38448 -6376 38468 -6368
rect 38476 -6376 38504 -6368
rect 38512 -6376 38532 -6368
rect 38688 -6368 38772 -6348
rect 38688 -6376 38708 -6368
rect 38716 -6376 38744 -6368
rect 38752 -6376 38772 -6368
rect 38808 -6368 38892 -6348
rect 38808 -6376 38828 -6368
rect 38836 -6376 38864 -6368
rect 38872 -6376 38892 -6368
rect 39048 -6368 39132 -6348
rect 39048 -6376 39068 -6368
rect 39076 -6376 39104 -6368
rect 39112 -6376 39132 -6368
rect 39168 -6368 39252 -6348
rect 39168 -6376 39188 -6368
rect 39196 -6376 39224 -6368
rect 39232 -6376 39252 -6368
rect 39408 -6368 39492 -6348
rect 39408 -6376 39428 -6368
rect 39436 -6376 39464 -6368
rect 39472 -6376 39492 -6368
rect 39528 -6368 39612 -6348
rect 39528 -6376 39548 -6368
rect 39556 -6376 39584 -6368
rect 39592 -6376 39612 -6368
rect 39768 -6368 39852 -6348
rect 39768 -6376 39788 -6368
rect 39796 -6376 39824 -6368
rect 39832 -6376 39852 -6368
rect 39888 -6368 39972 -6348
rect 39888 -6376 39908 -6368
rect 39916 -6376 39944 -6368
rect 39952 -6376 39972 -6368
rect 40128 -6368 40212 -6348
rect 40128 -6376 40148 -6368
rect 40156 -6376 40184 -6368
rect 40192 -6376 40212 -6368
rect 40248 -6368 40332 -6348
rect 40248 -6376 40268 -6368
rect 40276 -6376 40304 -6368
rect 40312 -6376 40332 -6368
rect 40488 -6368 40572 -6348
rect 40488 -6376 40508 -6368
rect 40516 -6376 40544 -6368
rect 40552 -6376 40572 -6368
rect 40608 -6368 40692 -6348
rect 40608 -6376 40628 -6368
rect 40636 -6376 40664 -6368
rect 40672 -6376 40692 -6368
rect 40848 -6368 40932 -6348
rect 40848 -6376 40868 -6368
rect 40876 -6376 40904 -6368
rect 40912 -6376 40932 -6368
rect 40968 -6368 41052 -6348
rect 40968 -6376 40988 -6368
rect 40996 -6376 41024 -6368
rect 41032 -6376 41052 -6368
rect 41208 -6368 41292 -6348
rect 41208 -6376 41228 -6368
rect 41236 -6376 41264 -6368
rect 41272 -6376 41292 -6368
rect 41328 -6368 41412 -6348
rect 41328 -6376 41348 -6368
rect 41356 -6376 41384 -6368
rect 41392 -6376 41412 -6368
rect 41568 -6368 41652 -6348
rect 41568 -6376 41588 -6368
rect 41596 -6376 41624 -6368
rect 41632 -6376 41652 -6368
rect 41688 -6368 41772 -6348
rect 41688 -6376 41708 -6368
rect 41716 -6376 41744 -6368
rect 41752 -6376 41772 -6368
rect 41928 -6368 42012 -6348
rect 41928 -6376 41948 -6368
rect 41956 -6376 41984 -6368
rect 41992 -6376 42012 -6368
rect 42048 -6368 42132 -6348
rect 42048 -6376 42068 -6368
rect 42076 -6376 42104 -6368
rect 42112 -6376 42132 -6368
rect 42288 -6368 42372 -6348
rect 42288 -6376 42308 -6368
rect 42316 -6376 42344 -6368
rect 42352 -6376 42372 -6368
rect 42408 -6368 42492 -6348
rect 42408 -6376 42428 -6368
rect 42436 -6376 42464 -6368
rect 42472 -6376 42492 -6368
rect 42648 -6368 42732 -6348
rect 42648 -6376 42668 -6368
rect 42676 -6376 42704 -6368
rect 42712 -6376 42732 -6368
rect 42768 -6368 42852 -6348
rect 42768 -6376 42788 -6368
rect 42796 -6376 42824 -6368
rect 42832 -6376 42852 -6368
rect 43008 -6368 43092 -6348
rect 43008 -6376 43028 -6368
rect 43036 -6376 43064 -6368
rect 43072 -6376 43092 -6368
rect 43128 -6368 43212 -6348
rect 43128 -6376 43148 -6368
rect 43156 -6376 43184 -6368
rect 43192 -6376 43212 -6368
rect 43248 -6368 43332 -6348
rect 43248 -6376 43268 -6368
rect 43276 -6376 43304 -6368
rect 43312 -6376 43332 -6368
rect 43488 -6368 43572 -6348
rect 43488 -6376 43508 -6368
rect 43516 -6376 43544 -6368
rect 43552 -6376 43572 -6368
rect 43608 -6368 43692 -6348
rect 43608 -6376 43628 -6368
rect 43636 -6376 43664 -6368
rect 43672 -6376 43692 -6368
rect 43848 -6368 43932 -6348
rect 43848 -6376 43868 -6368
rect 43876 -6376 43904 -6368
rect 43912 -6376 43932 -6368
rect 43968 -6368 44052 -6348
rect 43968 -6376 43988 -6368
rect 43996 -6376 44024 -6368
rect 44032 -6376 44052 -6368
rect 44208 -6368 44292 -6348
rect 44208 -6376 44228 -6368
rect 44236 -6376 44264 -6368
rect 44272 -6376 44292 -6368
rect 44328 -6368 44412 -6348
rect 44328 -6376 44348 -6368
rect 44356 -6376 44384 -6368
rect 44392 -6376 44412 -6368
rect 44448 -6368 44532 -6348
rect 44448 -6376 44468 -6368
rect 44476 -6376 44504 -6368
rect 44512 -6376 44532 -6368
rect 44688 -6368 44772 -6348
rect 44688 -6376 44708 -6368
rect 44716 -6376 44744 -6368
rect 44752 -6376 44772 -6368
rect 44808 -6368 44892 -6348
rect 44808 -6376 44828 -6368
rect 44836 -6376 44864 -6368
rect 44872 -6376 44892 -6368
rect 45048 -6368 45132 -6348
rect 45048 -6376 45068 -6368
rect 45076 -6376 45104 -6368
rect 45112 -6376 45132 -6368
rect 45168 -6368 45252 -6348
rect 45168 -6376 45188 -6368
rect 45196 -6376 45224 -6368
rect 45232 -6376 45252 -6368
rect 45408 -6368 45492 -6348
rect 45408 -6376 45428 -6368
rect 45436 -6376 45464 -6368
rect 45472 -6376 45492 -6368
rect 45528 -6368 45612 -6348
rect 45528 -6376 45548 -6368
rect 45556 -6376 45584 -6368
rect 45592 -6376 45612 -6368
rect 25876 -6404 25932 -6376
rect 26116 -6404 26172 -6376
rect 26236 -6404 26292 -6376
rect 26476 -6404 26532 -6376
rect 26596 -6404 26652 -6376
rect 26836 -6404 26892 -6376
rect 26956 -6404 27012 -6376
rect 27196 -6404 27252 -6376
rect 27316 -6404 27372 -6376
rect 27556 -6404 27612 -6376
rect 27676 -6404 27732 -6376
rect 27916 -6404 27972 -6376
rect 28036 -6404 28092 -6376
rect 28276 -6404 28332 -6376
rect 28396 -6404 28452 -6376
rect 28636 -6404 28692 -6376
rect 28756 -6404 28812 -6376
rect 28996 -6404 29052 -6376
rect 29116 -6404 29172 -6376
rect 29356 -6404 29412 -6376
rect 29476 -6404 29532 -6376
rect 29716 -6404 29772 -6376
rect 29836 -6404 29892 -6376
rect 30076 -6404 30132 -6376
rect 30196 -6404 30252 -6376
rect 30436 -6404 30492 -6376
rect 30556 -6404 30612 -6376
rect 30796 -6404 30852 -6376
rect 30916 -6404 30972 -6376
rect 31156 -6404 31212 -6376
rect 31276 -6404 31332 -6376
rect 31516 -6404 31572 -6376
rect 31636 -6404 31692 -6376
rect 31876 -6404 31932 -6376
rect 31996 -6404 32052 -6376
rect 32236 -6404 32292 -6376
rect 32356 -6404 32412 -6376
rect 32596 -6404 32652 -6376
rect 32716 -6404 32772 -6376
rect 32956 -6404 33012 -6376
rect 33076 -6404 33132 -6376
rect 33316 -6404 33372 -6376
rect 33436 -6404 33492 -6376
rect 33676 -6404 33732 -6376
rect 33796 -6404 33852 -6376
rect 34036 -6404 34092 -6376
rect 34156 -6404 34212 -6376
rect 34396 -6404 34452 -6376
rect 34516 -6404 34572 -6376
rect 34756 -6404 34812 -6376
rect 34876 -6404 34932 -6376
rect 35116 -6404 35172 -6376
rect 35236 -6404 35292 -6376
rect 35476 -6404 35532 -6376
rect 35596 -6404 35652 -6376
rect 35836 -6404 35892 -6376
rect 35956 -6404 36012 -6376
rect 36196 -6404 36252 -6376
rect 36316 -6404 36372 -6376
rect 36556 -6404 36612 -6376
rect 36676 -6404 36732 -6376
rect 36916 -6404 36972 -6376
rect 37036 -6404 37092 -6376
rect 37276 -6404 37332 -6376
rect 37396 -6404 37452 -6376
rect 37636 -6404 37692 -6376
rect 37756 -6404 37812 -6376
rect 37996 -6404 38052 -6376
rect 38116 -6404 38172 -6376
rect 38356 -6404 38412 -6376
rect 38476 -6404 38532 -6376
rect 38716 -6404 38772 -6376
rect 38836 -6404 38892 -6376
rect 39076 -6404 39132 -6376
rect 39196 -6404 39252 -6376
rect 39436 -6404 39492 -6376
rect 39556 -6404 39612 -6376
rect 39796 -6404 39852 -6376
rect 39916 -6404 39972 -6376
rect 40156 -6404 40212 -6376
rect 40276 -6404 40332 -6376
rect 40516 -6404 40572 -6376
rect 40636 -6404 40692 -6376
rect 40876 -6404 40932 -6376
rect 40996 -6404 41052 -6376
rect 41236 -6404 41292 -6376
rect 41356 -6404 41412 -6376
rect 41596 -6404 41652 -6376
rect 41716 -6404 41772 -6376
rect 41956 -6404 42012 -6376
rect 42076 -6404 42132 -6376
rect 42316 -6404 42372 -6376
rect 42436 -6404 42492 -6376
rect 42676 -6404 42732 -6376
rect 42796 -6404 42852 -6376
rect 43036 -6404 43092 -6376
rect 43156 -6404 43212 -6376
rect 43276 -6404 43332 -6376
rect 43516 -6404 43572 -6376
rect 43636 -6404 43692 -6376
rect 43876 -6404 43932 -6376
rect 43996 -6404 44052 -6376
rect 44236 -6404 44292 -6376
rect 44356 -6404 44412 -6376
rect 44476 -6404 44532 -6376
rect 44716 -6404 44772 -6376
rect 44836 -6404 44892 -6376
rect 45076 -6404 45132 -6376
rect 45196 -6404 45252 -6376
rect 45436 -6404 45492 -6376
rect 45556 -6404 45612 -6376
rect 25848 -6548 25932 -6528
rect 25848 -6556 25868 -6548
rect 25876 -6556 25904 -6548
rect 25912 -6556 25932 -6548
rect 25968 -6548 26052 -6528
rect 25968 -6556 25988 -6548
rect 25996 -6556 26024 -6548
rect 26032 -6556 26052 -6548
rect 26088 -6548 26172 -6528
rect 26088 -6556 26108 -6548
rect 26116 -6556 26144 -6548
rect 26152 -6556 26172 -6548
rect 26208 -6548 26292 -6528
rect 26208 -6556 26228 -6548
rect 26236 -6556 26264 -6548
rect 26272 -6556 26292 -6548
rect 26328 -6548 26412 -6528
rect 26328 -6556 26348 -6548
rect 26356 -6556 26384 -6548
rect 26392 -6556 26412 -6548
rect 26448 -6548 26532 -6528
rect 26448 -6556 26468 -6548
rect 26476 -6556 26504 -6548
rect 26512 -6556 26532 -6548
rect 26568 -6548 26652 -6528
rect 26568 -6556 26588 -6548
rect 26596 -6556 26624 -6548
rect 26632 -6556 26652 -6548
rect 26688 -6548 26772 -6528
rect 26688 -6556 26708 -6548
rect 26716 -6556 26744 -6548
rect 26752 -6556 26772 -6548
rect 26808 -6548 26892 -6528
rect 26808 -6556 26828 -6548
rect 26836 -6556 26864 -6548
rect 26872 -6556 26892 -6548
rect 26928 -6548 27012 -6528
rect 26928 -6556 26948 -6548
rect 26956 -6556 26984 -6548
rect 26992 -6556 27012 -6548
rect 27048 -6548 27132 -6528
rect 27048 -6556 27068 -6548
rect 27076 -6556 27104 -6548
rect 27112 -6556 27132 -6548
rect 27168 -6548 27252 -6528
rect 27168 -6556 27188 -6548
rect 27196 -6556 27224 -6548
rect 27232 -6556 27252 -6548
rect 27288 -6548 27372 -6528
rect 27288 -6556 27308 -6548
rect 27316 -6556 27344 -6548
rect 27352 -6556 27372 -6548
rect 27408 -6548 27492 -6528
rect 27408 -6556 27428 -6548
rect 27436 -6556 27464 -6548
rect 27472 -6556 27492 -6548
rect 27528 -6548 27612 -6528
rect 27528 -6556 27548 -6548
rect 27556 -6556 27584 -6548
rect 27592 -6556 27612 -6548
rect 27648 -6548 27732 -6528
rect 27648 -6556 27668 -6548
rect 27676 -6556 27704 -6548
rect 27712 -6556 27732 -6548
rect 27768 -6548 27852 -6528
rect 27768 -6556 27788 -6548
rect 27796 -6556 27824 -6548
rect 27832 -6556 27852 -6548
rect 27888 -6548 27972 -6528
rect 27888 -6556 27908 -6548
rect 27916 -6556 27944 -6548
rect 27952 -6556 27972 -6548
rect 28008 -6548 28092 -6528
rect 28008 -6556 28028 -6548
rect 28036 -6556 28064 -6548
rect 28072 -6556 28092 -6548
rect 28128 -6548 28212 -6528
rect 28128 -6556 28148 -6548
rect 28156 -6556 28184 -6548
rect 28192 -6556 28212 -6548
rect 28248 -6548 28332 -6528
rect 28248 -6556 28268 -6548
rect 28276 -6556 28304 -6548
rect 28312 -6556 28332 -6548
rect 28368 -6548 28452 -6528
rect 28368 -6556 28388 -6548
rect 28396 -6556 28424 -6548
rect 28432 -6556 28452 -6548
rect 28488 -6548 28572 -6528
rect 28488 -6556 28508 -6548
rect 28516 -6556 28544 -6548
rect 28552 -6556 28572 -6548
rect 28608 -6548 28692 -6528
rect 28608 -6556 28628 -6548
rect 28636 -6556 28664 -6548
rect 28672 -6556 28692 -6548
rect 28728 -6548 28812 -6528
rect 28728 -6556 28748 -6548
rect 28756 -6556 28784 -6548
rect 28792 -6556 28812 -6548
rect 28848 -6548 28932 -6528
rect 28848 -6556 28868 -6548
rect 28876 -6556 28904 -6548
rect 28912 -6556 28932 -6548
rect 28968 -6548 29052 -6528
rect 28968 -6556 28988 -6548
rect 28996 -6556 29024 -6548
rect 29032 -6556 29052 -6548
rect 29088 -6548 29172 -6528
rect 29088 -6556 29108 -6548
rect 29116 -6556 29144 -6548
rect 29152 -6556 29172 -6548
rect 29208 -6548 29292 -6528
rect 29208 -6556 29228 -6548
rect 29236 -6556 29264 -6548
rect 29272 -6556 29292 -6548
rect 29328 -6548 29412 -6528
rect 29328 -6556 29348 -6548
rect 29356 -6556 29384 -6548
rect 29392 -6556 29412 -6548
rect 29448 -6548 29532 -6528
rect 29448 -6556 29468 -6548
rect 29476 -6556 29504 -6548
rect 29512 -6556 29532 -6548
rect 29568 -6548 29652 -6528
rect 29568 -6556 29588 -6548
rect 29596 -6556 29624 -6548
rect 29632 -6556 29652 -6548
rect 29688 -6548 29772 -6528
rect 29688 -6556 29708 -6548
rect 29716 -6556 29744 -6548
rect 29752 -6556 29772 -6548
rect 29808 -6548 29892 -6528
rect 29808 -6556 29828 -6548
rect 29836 -6556 29864 -6548
rect 29872 -6556 29892 -6548
rect 29928 -6548 30012 -6528
rect 29928 -6556 29948 -6548
rect 29956 -6556 29984 -6548
rect 29992 -6556 30012 -6548
rect 30048 -6548 30132 -6528
rect 30048 -6556 30068 -6548
rect 30076 -6556 30104 -6548
rect 30112 -6556 30132 -6548
rect 30168 -6548 30252 -6528
rect 30168 -6556 30188 -6548
rect 30196 -6556 30224 -6548
rect 30232 -6556 30252 -6548
rect 30288 -6548 30372 -6528
rect 30288 -6556 30308 -6548
rect 30316 -6556 30344 -6548
rect 30352 -6556 30372 -6548
rect 30408 -6548 30492 -6528
rect 30408 -6556 30428 -6548
rect 30436 -6556 30464 -6548
rect 30472 -6556 30492 -6548
rect 30528 -6548 30612 -6528
rect 30528 -6556 30548 -6548
rect 30556 -6556 30584 -6548
rect 30592 -6556 30612 -6548
rect 30648 -6548 30732 -6528
rect 30648 -6556 30668 -6548
rect 30676 -6556 30704 -6548
rect 30712 -6556 30732 -6548
rect 30768 -6548 30852 -6528
rect 30768 -6556 30788 -6548
rect 30796 -6556 30824 -6548
rect 30832 -6556 30852 -6548
rect 30888 -6548 30972 -6528
rect 30888 -6556 30908 -6548
rect 30916 -6556 30944 -6548
rect 30952 -6556 30972 -6548
rect 31008 -6548 31092 -6528
rect 31008 -6556 31028 -6548
rect 31036 -6556 31064 -6548
rect 31072 -6556 31092 -6548
rect 31128 -6548 31212 -6528
rect 31128 -6556 31148 -6548
rect 31156 -6556 31184 -6548
rect 31192 -6556 31212 -6548
rect 31248 -6548 31332 -6528
rect 31248 -6556 31268 -6548
rect 31276 -6556 31304 -6548
rect 31312 -6556 31332 -6548
rect 31368 -6548 31452 -6528
rect 31368 -6556 31388 -6548
rect 31396 -6556 31424 -6548
rect 31432 -6556 31452 -6548
rect 31488 -6548 31572 -6528
rect 31488 -6556 31508 -6548
rect 31516 -6556 31544 -6548
rect 31552 -6556 31572 -6548
rect 31608 -6548 31692 -6528
rect 31608 -6556 31628 -6548
rect 31636 -6556 31664 -6548
rect 31672 -6556 31692 -6548
rect 31728 -6548 31812 -6528
rect 31728 -6556 31748 -6548
rect 31756 -6556 31784 -6548
rect 31792 -6556 31812 -6548
rect 31848 -6548 31932 -6528
rect 31848 -6556 31868 -6548
rect 31876 -6556 31904 -6548
rect 31912 -6556 31932 -6548
rect 31968 -6548 32052 -6528
rect 31968 -6556 31988 -6548
rect 31996 -6556 32024 -6548
rect 32032 -6556 32052 -6548
rect 32088 -6548 32172 -6528
rect 32088 -6556 32108 -6548
rect 32116 -6556 32144 -6548
rect 32152 -6556 32172 -6548
rect 32208 -6548 32292 -6528
rect 32208 -6556 32228 -6548
rect 32236 -6556 32264 -6548
rect 32272 -6556 32292 -6548
rect 32328 -6548 32412 -6528
rect 32328 -6556 32348 -6548
rect 32356 -6556 32384 -6548
rect 32392 -6556 32412 -6548
rect 32448 -6548 32532 -6528
rect 32448 -6556 32468 -6548
rect 32476 -6556 32504 -6548
rect 32512 -6556 32532 -6548
rect 32568 -6548 32652 -6528
rect 32568 -6556 32588 -6548
rect 32596 -6556 32624 -6548
rect 32632 -6556 32652 -6548
rect 32688 -6548 32772 -6528
rect 32688 -6556 32708 -6548
rect 32716 -6556 32744 -6548
rect 32752 -6556 32772 -6548
rect 32808 -6548 32892 -6528
rect 32808 -6556 32828 -6548
rect 32836 -6556 32864 -6548
rect 32872 -6556 32892 -6548
rect 32928 -6548 33012 -6528
rect 32928 -6556 32948 -6548
rect 32956 -6556 32984 -6548
rect 32992 -6556 33012 -6548
rect 33048 -6548 33132 -6528
rect 33048 -6556 33068 -6548
rect 33076 -6556 33104 -6548
rect 33112 -6556 33132 -6548
rect 33168 -6548 33252 -6528
rect 33168 -6556 33188 -6548
rect 33196 -6556 33224 -6548
rect 33232 -6556 33252 -6548
rect 33288 -6548 33372 -6528
rect 33288 -6556 33308 -6548
rect 33316 -6556 33344 -6548
rect 33352 -6556 33372 -6548
rect 33408 -6548 33492 -6528
rect 33408 -6556 33428 -6548
rect 33436 -6556 33464 -6548
rect 33472 -6556 33492 -6548
rect 33528 -6548 33612 -6528
rect 33528 -6556 33548 -6548
rect 33556 -6556 33584 -6548
rect 33592 -6556 33612 -6548
rect 33648 -6548 33732 -6528
rect 33648 -6556 33668 -6548
rect 33676 -6556 33704 -6548
rect 33712 -6556 33732 -6548
rect 33768 -6548 33852 -6528
rect 33768 -6556 33788 -6548
rect 33796 -6556 33824 -6548
rect 33832 -6556 33852 -6548
rect 33888 -6548 33972 -6528
rect 33888 -6556 33908 -6548
rect 33916 -6556 33944 -6548
rect 33952 -6556 33972 -6548
rect 34008 -6548 34092 -6528
rect 34008 -6556 34028 -6548
rect 34036 -6556 34064 -6548
rect 34072 -6556 34092 -6548
rect 34128 -6548 34212 -6528
rect 34128 -6556 34148 -6548
rect 34156 -6556 34184 -6548
rect 34192 -6556 34212 -6548
rect 34248 -6548 34332 -6528
rect 34248 -6556 34268 -6548
rect 34276 -6556 34304 -6548
rect 34312 -6556 34332 -6548
rect 34368 -6548 34452 -6528
rect 34368 -6556 34388 -6548
rect 34396 -6556 34424 -6548
rect 34432 -6556 34452 -6548
rect 34488 -6548 34572 -6528
rect 34488 -6556 34508 -6548
rect 34516 -6556 34544 -6548
rect 34552 -6556 34572 -6548
rect 34608 -6548 34692 -6528
rect 34608 -6556 34628 -6548
rect 34636 -6556 34664 -6548
rect 34672 -6556 34692 -6548
rect 34728 -6548 34812 -6528
rect 34728 -6556 34748 -6548
rect 34756 -6556 34784 -6548
rect 34792 -6556 34812 -6548
rect 34848 -6548 34932 -6528
rect 34848 -6556 34868 -6548
rect 34876 -6556 34904 -6548
rect 34912 -6556 34932 -6548
rect 34968 -6548 35052 -6528
rect 34968 -6556 34988 -6548
rect 34996 -6556 35024 -6548
rect 35032 -6556 35052 -6548
rect 35088 -6548 35172 -6528
rect 35088 -6556 35108 -6548
rect 35116 -6556 35144 -6548
rect 35152 -6556 35172 -6548
rect 35208 -6548 35292 -6528
rect 35208 -6556 35228 -6548
rect 35236 -6556 35264 -6548
rect 35272 -6556 35292 -6548
rect 35328 -6548 35412 -6528
rect 35328 -6556 35348 -6548
rect 35356 -6556 35384 -6548
rect 35392 -6556 35412 -6548
rect 35448 -6548 35532 -6528
rect 35448 -6556 35468 -6548
rect 35476 -6556 35504 -6548
rect 35512 -6556 35532 -6548
rect 35568 -6548 35652 -6528
rect 35568 -6556 35588 -6548
rect 35596 -6556 35624 -6548
rect 35632 -6556 35652 -6548
rect 35688 -6548 35772 -6528
rect 35688 -6556 35708 -6548
rect 35716 -6556 35744 -6548
rect 35752 -6556 35772 -6548
rect 35808 -6548 35892 -6528
rect 35808 -6556 35828 -6548
rect 35836 -6556 35864 -6548
rect 35872 -6556 35892 -6548
rect 35928 -6548 36012 -6528
rect 35928 -6556 35948 -6548
rect 35956 -6556 35984 -6548
rect 35992 -6556 36012 -6548
rect 36048 -6548 36132 -6528
rect 36048 -6556 36068 -6548
rect 36076 -6556 36104 -6548
rect 36112 -6556 36132 -6548
rect 36168 -6548 36252 -6528
rect 36168 -6556 36188 -6548
rect 36196 -6556 36224 -6548
rect 36232 -6556 36252 -6548
rect 36288 -6548 36372 -6528
rect 36288 -6556 36308 -6548
rect 36316 -6556 36344 -6548
rect 36352 -6556 36372 -6548
rect 36408 -6548 36492 -6528
rect 36408 -6556 36428 -6548
rect 36436 -6556 36464 -6548
rect 36472 -6556 36492 -6548
rect 36528 -6548 36612 -6528
rect 36528 -6556 36548 -6548
rect 36556 -6556 36584 -6548
rect 36592 -6556 36612 -6548
rect 36648 -6548 36732 -6528
rect 36648 -6556 36668 -6548
rect 36676 -6556 36704 -6548
rect 36712 -6556 36732 -6548
rect 36768 -6548 36852 -6528
rect 36768 -6556 36788 -6548
rect 36796 -6556 36824 -6548
rect 36832 -6556 36852 -6548
rect 36888 -6548 36972 -6528
rect 36888 -6556 36908 -6548
rect 36916 -6556 36944 -6548
rect 36952 -6556 36972 -6548
rect 37008 -6548 37092 -6528
rect 37008 -6556 37028 -6548
rect 37036 -6556 37064 -6548
rect 37072 -6556 37092 -6548
rect 37128 -6548 37212 -6528
rect 37128 -6556 37148 -6548
rect 37156 -6556 37184 -6548
rect 37192 -6556 37212 -6548
rect 37248 -6548 37332 -6528
rect 37248 -6556 37268 -6548
rect 37276 -6556 37304 -6548
rect 37312 -6556 37332 -6548
rect 37368 -6548 37452 -6528
rect 37368 -6556 37388 -6548
rect 37396 -6556 37424 -6548
rect 37432 -6556 37452 -6548
rect 37488 -6548 37572 -6528
rect 37488 -6556 37508 -6548
rect 37516 -6556 37544 -6548
rect 37552 -6556 37572 -6548
rect 37608 -6548 37692 -6528
rect 37608 -6556 37628 -6548
rect 37636 -6556 37664 -6548
rect 37672 -6556 37692 -6548
rect 37728 -6548 37812 -6528
rect 37728 -6556 37748 -6548
rect 37756 -6556 37784 -6548
rect 37792 -6556 37812 -6548
rect 37848 -6548 37932 -6528
rect 37848 -6556 37868 -6548
rect 37876 -6556 37904 -6548
rect 37912 -6556 37932 -6548
rect 37968 -6548 38052 -6528
rect 37968 -6556 37988 -6548
rect 37996 -6556 38024 -6548
rect 38032 -6556 38052 -6548
rect 38088 -6548 38172 -6528
rect 38088 -6556 38108 -6548
rect 38116 -6556 38144 -6548
rect 38152 -6556 38172 -6548
rect 38208 -6548 38292 -6528
rect 38208 -6556 38228 -6548
rect 38236 -6556 38264 -6548
rect 38272 -6556 38292 -6548
rect 38328 -6548 38412 -6528
rect 38328 -6556 38348 -6548
rect 38356 -6556 38384 -6548
rect 38392 -6556 38412 -6548
rect 38448 -6548 38532 -6528
rect 38448 -6556 38468 -6548
rect 38476 -6556 38504 -6548
rect 38512 -6556 38532 -6548
rect 38568 -6548 38652 -6528
rect 38568 -6556 38588 -6548
rect 38596 -6556 38624 -6548
rect 38632 -6556 38652 -6548
rect 38688 -6548 38772 -6528
rect 38688 -6556 38708 -6548
rect 38716 -6556 38744 -6548
rect 38752 -6556 38772 -6548
rect 38808 -6548 38892 -6528
rect 38808 -6556 38828 -6548
rect 38836 -6556 38864 -6548
rect 38872 -6556 38892 -6548
rect 38928 -6548 39012 -6528
rect 38928 -6556 38948 -6548
rect 38956 -6556 38984 -6548
rect 38992 -6556 39012 -6548
rect 39048 -6548 39132 -6528
rect 39048 -6556 39068 -6548
rect 39076 -6556 39104 -6548
rect 39112 -6556 39132 -6548
rect 39168 -6548 39252 -6528
rect 39168 -6556 39188 -6548
rect 39196 -6556 39224 -6548
rect 39232 -6556 39252 -6548
rect 39288 -6548 39372 -6528
rect 39288 -6556 39308 -6548
rect 39316 -6556 39344 -6548
rect 39352 -6556 39372 -6548
rect 39408 -6548 39492 -6528
rect 39408 -6556 39428 -6548
rect 39436 -6556 39464 -6548
rect 39472 -6556 39492 -6548
rect 39528 -6548 39612 -6528
rect 39528 -6556 39548 -6548
rect 39556 -6556 39584 -6548
rect 39592 -6556 39612 -6548
rect 39648 -6548 39732 -6528
rect 39648 -6556 39668 -6548
rect 39676 -6556 39704 -6548
rect 39712 -6556 39732 -6548
rect 39768 -6548 39852 -6528
rect 39768 -6556 39788 -6548
rect 39796 -6556 39824 -6548
rect 39832 -6556 39852 -6548
rect 39888 -6548 39972 -6528
rect 39888 -6556 39908 -6548
rect 39916 -6556 39944 -6548
rect 39952 -6556 39972 -6548
rect 40008 -6548 40092 -6528
rect 40008 -6556 40028 -6548
rect 40036 -6556 40064 -6548
rect 40072 -6556 40092 -6548
rect 40128 -6548 40212 -6528
rect 40128 -6556 40148 -6548
rect 40156 -6556 40184 -6548
rect 40192 -6556 40212 -6548
rect 40248 -6548 40332 -6528
rect 40248 -6556 40268 -6548
rect 40276 -6556 40304 -6548
rect 40312 -6556 40332 -6548
rect 40368 -6548 40452 -6528
rect 40368 -6556 40388 -6548
rect 40396 -6556 40424 -6548
rect 40432 -6556 40452 -6548
rect 40488 -6548 40572 -6528
rect 40488 -6556 40508 -6548
rect 40516 -6556 40544 -6548
rect 40552 -6556 40572 -6548
rect 40608 -6548 40692 -6528
rect 40608 -6556 40628 -6548
rect 40636 -6556 40664 -6548
rect 40672 -6556 40692 -6548
rect 40728 -6548 40812 -6528
rect 40728 -6556 40748 -6548
rect 40756 -6556 40784 -6548
rect 40792 -6556 40812 -6548
rect 40848 -6548 40932 -6528
rect 40848 -6556 40868 -6548
rect 40876 -6556 40904 -6548
rect 40912 -6556 40932 -6548
rect 40968 -6548 41052 -6528
rect 40968 -6556 40988 -6548
rect 40996 -6556 41024 -6548
rect 41032 -6556 41052 -6548
rect 41088 -6548 41172 -6528
rect 41088 -6556 41108 -6548
rect 41116 -6556 41144 -6548
rect 41152 -6556 41172 -6548
rect 41208 -6548 41292 -6528
rect 41208 -6556 41228 -6548
rect 41236 -6556 41264 -6548
rect 41272 -6556 41292 -6548
rect 41328 -6548 41412 -6528
rect 41328 -6556 41348 -6548
rect 41356 -6556 41384 -6548
rect 41392 -6556 41412 -6548
rect 41448 -6548 41532 -6528
rect 41448 -6556 41468 -6548
rect 41476 -6556 41504 -6548
rect 41512 -6556 41532 -6548
rect 41568 -6548 41652 -6528
rect 41568 -6556 41588 -6548
rect 41596 -6556 41624 -6548
rect 41632 -6556 41652 -6548
rect 41688 -6548 41772 -6528
rect 41688 -6556 41708 -6548
rect 41716 -6556 41744 -6548
rect 41752 -6556 41772 -6548
rect 41808 -6548 41892 -6528
rect 41808 -6556 41828 -6548
rect 41836 -6556 41864 -6548
rect 41872 -6556 41892 -6548
rect 41928 -6548 42012 -6528
rect 41928 -6556 41948 -6548
rect 41956 -6556 41984 -6548
rect 41992 -6556 42012 -6548
rect 42048 -6548 42132 -6528
rect 42048 -6556 42068 -6548
rect 42076 -6556 42104 -6548
rect 42112 -6556 42132 -6548
rect 42168 -6548 42252 -6528
rect 42168 -6556 42188 -6548
rect 42196 -6556 42224 -6548
rect 42232 -6556 42252 -6548
rect 42288 -6548 42372 -6528
rect 42288 -6556 42308 -6548
rect 42316 -6556 42344 -6548
rect 42352 -6556 42372 -6548
rect 42408 -6548 42492 -6528
rect 42408 -6556 42428 -6548
rect 42436 -6556 42464 -6548
rect 42472 -6556 42492 -6548
rect 42528 -6548 42612 -6528
rect 42528 -6556 42548 -6548
rect 42556 -6556 42584 -6548
rect 42592 -6556 42612 -6548
rect 42648 -6548 42732 -6528
rect 42648 -6556 42668 -6548
rect 42676 -6556 42704 -6548
rect 42712 -6556 42732 -6548
rect 42768 -6548 42852 -6528
rect 42768 -6556 42788 -6548
rect 42796 -6556 42824 -6548
rect 42832 -6556 42852 -6548
rect 42888 -6548 42972 -6528
rect 42888 -6556 42908 -6548
rect 42916 -6556 42944 -6548
rect 42952 -6556 42972 -6548
rect 43008 -6548 43092 -6528
rect 43008 -6556 43028 -6548
rect 43036 -6556 43064 -6548
rect 43072 -6556 43092 -6548
rect 43128 -6548 43212 -6528
rect 43128 -6556 43148 -6548
rect 43156 -6556 43184 -6548
rect 43192 -6556 43212 -6548
rect 43248 -6548 43332 -6528
rect 43248 -6556 43268 -6548
rect 43276 -6556 43304 -6548
rect 43312 -6556 43332 -6548
rect 43368 -6548 43452 -6528
rect 43368 -6556 43388 -6548
rect 43396 -6556 43424 -6548
rect 43432 -6556 43452 -6548
rect 43488 -6548 43572 -6528
rect 43488 -6556 43508 -6548
rect 43516 -6556 43544 -6548
rect 43552 -6556 43572 -6548
rect 43608 -6548 43692 -6528
rect 43608 -6556 43628 -6548
rect 43636 -6556 43664 -6548
rect 43672 -6556 43692 -6548
rect 43728 -6548 43812 -6528
rect 43728 -6556 43748 -6548
rect 43756 -6556 43784 -6548
rect 43792 -6556 43812 -6548
rect 43848 -6548 43932 -6528
rect 43848 -6556 43868 -6548
rect 43876 -6556 43904 -6548
rect 43912 -6556 43932 -6548
rect 43968 -6548 44052 -6528
rect 43968 -6556 43988 -6548
rect 43996 -6556 44024 -6548
rect 44032 -6556 44052 -6548
rect 44088 -6548 44172 -6528
rect 44088 -6556 44108 -6548
rect 44116 -6556 44144 -6548
rect 44152 -6556 44172 -6548
rect 44208 -6548 44292 -6528
rect 44208 -6556 44228 -6548
rect 44236 -6556 44264 -6548
rect 44272 -6556 44292 -6548
rect 44328 -6548 44412 -6528
rect 44328 -6556 44348 -6548
rect 44356 -6556 44384 -6548
rect 44392 -6556 44412 -6548
rect 44448 -6548 44532 -6528
rect 44448 -6556 44468 -6548
rect 44476 -6556 44504 -6548
rect 44512 -6556 44532 -6548
rect 44568 -6548 44652 -6528
rect 44568 -6556 44588 -6548
rect 44596 -6556 44624 -6548
rect 44632 -6556 44652 -6548
rect 44688 -6548 44772 -6528
rect 44688 -6556 44708 -6548
rect 44716 -6556 44744 -6548
rect 44752 -6556 44772 -6548
rect 44808 -6548 44892 -6528
rect 44808 -6556 44828 -6548
rect 44836 -6556 44864 -6548
rect 44872 -6556 44892 -6548
rect 44928 -6548 45012 -6528
rect 44928 -6556 44948 -6548
rect 44956 -6556 44984 -6548
rect 44992 -6556 45012 -6548
rect 45048 -6548 45132 -6528
rect 45048 -6556 45068 -6548
rect 45076 -6556 45104 -6548
rect 45112 -6556 45132 -6548
rect 45168 -6548 45252 -6528
rect 45168 -6556 45188 -6548
rect 45196 -6556 45224 -6548
rect 45232 -6556 45252 -6548
rect 45288 -6548 45372 -6528
rect 45288 -6556 45308 -6548
rect 45316 -6556 45344 -6548
rect 45352 -6556 45372 -6548
rect 45408 -6548 45492 -6528
rect 45408 -6556 45428 -6548
rect 45436 -6556 45464 -6548
rect 45472 -6556 45492 -6548
rect 45528 -6548 45612 -6528
rect 45528 -6556 45548 -6548
rect 45556 -6556 45584 -6548
rect 45592 -6556 45612 -6548
rect 25876 -6584 25932 -6556
rect 25996 -6584 26052 -6556
rect 26116 -6584 26172 -6556
rect 26236 -6584 26292 -6556
rect 26356 -6584 26412 -6556
rect 26476 -6584 26532 -6556
rect 26596 -6584 26652 -6556
rect 26716 -6584 26772 -6556
rect 26836 -6584 26892 -6556
rect 26956 -6584 27012 -6556
rect 27076 -6584 27132 -6556
rect 27196 -6584 27252 -6556
rect 27316 -6584 27372 -6556
rect 27436 -6584 27492 -6556
rect 27556 -6584 27612 -6556
rect 27676 -6584 27732 -6556
rect 27796 -6584 27852 -6556
rect 27916 -6584 27972 -6556
rect 28036 -6584 28092 -6556
rect 28156 -6584 28212 -6556
rect 28276 -6584 28332 -6556
rect 28396 -6584 28452 -6556
rect 28516 -6584 28572 -6556
rect 28636 -6584 28692 -6556
rect 28756 -6584 28812 -6556
rect 28876 -6584 28932 -6556
rect 28996 -6584 29052 -6556
rect 29116 -6584 29172 -6556
rect 29236 -6584 29292 -6556
rect 29356 -6584 29412 -6556
rect 29476 -6584 29532 -6556
rect 29596 -6584 29652 -6556
rect 29716 -6584 29772 -6556
rect 29836 -6584 29892 -6556
rect 29956 -6584 30012 -6556
rect 30076 -6584 30132 -6556
rect 30196 -6584 30252 -6556
rect 30316 -6584 30372 -6556
rect 30436 -6584 30492 -6556
rect 30556 -6584 30612 -6556
rect 30676 -6584 30732 -6556
rect 30796 -6584 30852 -6556
rect 30916 -6584 30972 -6556
rect 31036 -6584 31092 -6556
rect 31156 -6584 31212 -6556
rect 31276 -6584 31332 -6556
rect 31396 -6584 31452 -6556
rect 31516 -6584 31572 -6556
rect 31636 -6584 31692 -6556
rect 31756 -6584 31812 -6556
rect 31876 -6584 31932 -6556
rect 31996 -6584 32052 -6556
rect 32116 -6584 32172 -6556
rect 32236 -6584 32292 -6556
rect 32356 -6584 32412 -6556
rect 32476 -6584 32532 -6556
rect 32596 -6584 32652 -6556
rect 32716 -6584 32772 -6556
rect 32836 -6584 32892 -6556
rect 32956 -6584 33012 -6556
rect 33076 -6584 33132 -6556
rect 33196 -6584 33252 -6556
rect 33316 -6584 33372 -6556
rect 33436 -6584 33492 -6556
rect 33556 -6584 33612 -6556
rect 33676 -6584 33732 -6556
rect 33796 -6584 33852 -6556
rect 33916 -6584 33972 -6556
rect 34036 -6584 34092 -6556
rect 34156 -6584 34212 -6556
rect 34276 -6584 34332 -6556
rect 34396 -6584 34452 -6556
rect 34516 -6584 34572 -6556
rect 34636 -6584 34692 -6556
rect 34756 -6584 34812 -6556
rect 34876 -6584 34932 -6556
rect 34996 -6584 35052 -6556
rect 35116 -6584 35172 -6556
rect 35236 -6584 35292 -6556
rect 35356 -6584 35412 -6556
rect 35476 -6584 35532 -6556
rect 35596 -6584 35652 -6556
rect 35716 -6584 35772 -6556
rect 35836 -6584 35892 -6556
rect 35956 -6584 36012 -6556
rect 36076 -6584 36132 -6556
rect 36196 -6584 36252 -6556
rect 36316 -6584 36372 -6556
rect 36436 -6584 36492 -6556
rect 36556 -6584 36612 -6556
rect 36676 -6584 36732 -6556
rect 36796 -6584 36852 -6556
rect 36916 -6584 36972 -6556
rect 37036 -6584 37092 -6556
rect 37156 -6584 37212 -6556
rect 37276 -6584 37332 -6556
rect 37396 -6584 37452 -6556
rect 37516 -6584 37572 -6556
rect 37636 -6584 37692 -6556
rect 37756 -6584 37812 -6556
rect 37876 -6584 37932 -6556
rect 37996 -6584 38052 -6556
rect 38116 -6584 38172 -6556
rect 38236 -6584 38292 -6556
rect 38356 -6584 38412 -6556
rect 38476 -6584 38532 -6556
rect 38596 -6584 38652 -6556
rect 38716 -6584 38772 -6556
rect 38836 -6584 38892 -6556
rect 38956 -6584 39012 -6556
rect 39076 -6584 39132 -6556
rect 39196 -6584 39252 -6556
rect 39316 -6584 39372 -6556
rect 39436 -6584 39492 -6556
rect 39556 -6584 39612 -6556
rect 39676 -6584 39732 -6556
rect 39796 -6584 39852 -6556
rect 39916 -6584 39972 -6556
rect 40036 -6584 40092 -6556
rect 40156 -6584 40212 -6556
rect 40276 -6584 40332 -6556
rect 40396 -6584 40452 -6556
rect 40516 -6584 40572 -6556
rect 40636 -6584 40692 -6556
rect 40756 -6584 40812 -6556
rect 40876 -6584 40932 -6556
rect 40996 -6584 41052 -6556
rect 41116 -6584 41172 -6556
rect 41236 -6584 41292 -6556
rect 41356 -6584 41412 -6556
rect 41476 -6584 41532 -6556
rect 41596 -6584 41652 -6556
rect 41716 -6584 41772 -6556
rect 41836 -6584 41892 -6556
rect 41956 -6584 42012 -6556
rect 42076 -6584 42132 -6556
rect 42196 -6584 42252 -6556
rect 42316 -6584 42372 -6556
rect 42436 -6584 42492 -6556
rect 42556 -6584 42612 -6556
rect 42676 -6584 42732 -6556
rect 42796 -6584 42852 -6556
rect 42916 -6584 42972 -6556
rect 43036 -6584 43092 -6556
rect 43156 -6584 43212 -6556
rect 43276 -6584 43332 -6556
rect 43396 -6584 43452 -6556
rect 43516 -6584 43572 -6556
rect 43636 -6584 43692 -6556
rect 43756 -6584 43812 -6556
rect 43876 -6584 43932 -6556
rect 43996 -6584 44052 -6556
rect 44116 -6584 44172 -6556
rect 44236 -6584 44292 -6556
rect 44356 -6584 44412 -6556
rect 44476 -6584 44532 -6556
rect 44596 -6584 44652 -6556
rect 44716 -6584 44772 -6556
rect 44836 -6584 44892 -6556
rect 44956 -6584 45012 -6556
rect 45076 -6584 45132 -6556
rect 45196 -6584 45252 -6556
rect 45316 -6584 45372 -6556
rect 45436 -6584 45492 -6556
rect 45556 -6584 45612 -6556
rect 25848 -6728 25932 -6708
rect 25848 -6736 25868 -6728
rect 25876 -6736 25904 -6728
rect 25912 -6736 25932 -6728
rect 25968 -6728 26052 -6708
rect 25968 -6736 25988 -6728
rect 25996 -6736 26024 -6728
rect 26032 -6736 26052 -6728
rect 26088 -6728 26172 -6708
rect 26088 -6736 26108 -6728
rect 26116 -6736 26144 -6728
rect 26152 -6736 26172 -6728
rect 26208 -6728 26292 -6708
rect 26208 -6736 26228 -6728
rect 26236 -6736 26264 -6728
rect 26272 -6736 26292 -6728
rect 26328 -6728 26412 -6708
rect 26328 -6736 26348 -6728
rect 26356 -6736 26384 -6728
rect 26392 -6736 26412 -6728
rect 26448 -6728 26532 -6708
rect 26448 -6736 26468 -6728
rect 26476 -6736 26504 -6728
rect 26512 -6736 26532 -6728
rect 26568 -6728 26652 -6708
rect 26568 -6736 26588 -6728
rect 26596 -6736 26624 -6728
rect 26632 -6736 26652 -6728
rect 26688 -6728 26772 -6708
rect 26688 -6736 26708 -6728
rect 26716 -6736 26744 -6728
rect 26752 -6736 26772 -6728
rect 26808 -6728 26892 -6708
rect 26808 -6736 26828 -6728
rect 26836 -6736 26864 -6728
rect 26872 -6736 26892 -6728
rect 26928 -6728 27012 -6708
rect 26928 -6736 26948 -6728
rect 26956 -6736 26984 -6728
rect 26992 -6736 27012 -6728
rect 27048 -6728 27132 -6708
rect 27048 -6736 27068 -6728
rect 27076 -6736 27104 -6728
rect 27112 -6736 27132 -6728
rect 27168 -6728 27252 -6708
rect 27168 -6736 27188 -6728
rect 27196 -6736 27224 -6728
rect 27232 -6736 27252 -6728
rect 27288 -6728 27372 -6708
rect 27288 -6736 27308 -6728
rect 27316 -6736 27344 -6728
rect 27352 -6736 27372 -6728
rect 27408 -6728 27492 -6708
rect 27408 -6736 27428 -6728
rect 27436 -6736 27464 -6728
rect 27472 -6736 27492 -6728
rect 27528 -6728 27612 -6708
rect 27528 -6736 27548 -6728
rect 27556 -6736 27584 -6728
rect 27592 -6736 27612 -6728
rect 27648 -6728 27732 -6708
rect 27648 -6736 27668 -6728
rect 27676 -6736 27704 -6728
rect 27712 -6736 27732 -6728
rect 27768 -6728 27852 -6708
rect 27768 -6736 27788 -6728
rect 27796 -6736 27824 -6728
rect 27832 -6736 27852 -6728
rect 27888 -6728 27972 -6708
rect 27888 -6736 27908 -6728
rect 27916 -6736 27944 -6728
rect 27952 -6736 27972 -6728
rect 28008 -6728 28092 -6708
rect 28008 -6736 28028 -6728
rect 28036 -6736 28064 -6728
rect 28072 -6736 28092 -6728
rect 28128 -6728 28212 -6708
rect 28128 -6736 28148 -6728
rect 28156 -6736 28184 -6728
rect 28192 -6736 28212 -6728
rect 28248 -6728 28332 -6708
rect 28248 -6736 28268 -6728
rect 28276 -6736 28304 -6728
rect 28312 -6736 28332 -6728
rect 28368 -6728 28452 -6708
rect 28368 -6736 28388 -6728
rect 28396 -6736 28424 -6728
rect 28432 -6736 28452 -6728
rect 28488 -6728 28572 -6708
rect 28488 -6736 28508 -6728
rect 28516 -6736 28544 -6728
rect 28552 -6736 28572 -6728
rect 28608 -6728 28692 -6708
rect 28608 -6736 28628 -6728
rect 28636 -6736 28664 -6728
rect 28672 -6736 28692 -6728
rect 28728 -6728 28812 -6708
rect 28728 -6736 28748 -6728
rect 28756 -6736 28784 -6728
rect 28792 -6736 28812 -6728
rect 28848 -6728 28932 -6708
rect 28848 -6736 28868 -6728
rect 28876 -6736 28904 -6728
rect 28912 -6736 28932 -6728
rect 28968 -6728 29052 -6708
rect 28968 -6736 28988 -6728
rect 28996 -6736 29024 -6728
rect 29032 -6736 29052 -6728
rect 29088 -6728 29172 -6708
rect 29088 -6736 29108 -6728
rect 29116 -6736 29144 -6728
rect 29152 -6736 29172 -6728
rect 29208 -6728 29292 -6708
rect 29208 -6736 29228 -6728
rect 29236 -6736 29264 -6728
rect 29272 -6736 29292 -6728
rect 29328 -6728 29412 -6708
rect 29328 -6736 29348 -6728
rect 29356 -6736 29384 -6728
rect 29392 -6736 29412 -6728
rect 29448 -6728 29532 -6708
rect 29448 -6736 29468 -6728
rect 29476 -6736 29504 -6728
rect 29512 -6736 29532 -6728
rect 29568 -6728 29652 -6708
rect 29568 -6736 29588 -6728
rect 29596 -6736 29624 -6728
rect 29632 -6736 29652 -6728
rect 29688 -6728 29772 -6708
rect 29688 -6736 29708 -6728
rect 29716 -6736 29744 -6728
rect 29752 -6736 29772 -6728
rect 29808 -6728 29892 -6708
rect 29808 -6736 29828 -6728
rect 29836 -6736 29864 -6728
rect 29872 -6736 29892 -6728
rect 29928 -6728 30012 -6708
rect 29928 -6736 29948 -6728
rect 29956 -6736 29984 -6728
rect 29992 -6736 30012 -6728
rect 30048 -6728 30132 -6708
rect 30048 -6736 30068 -6728
rect 30076 -6736 30104 -6728
rect 30112 -6736 30132 -6728
rect 30168 -6728 30252 -6708
rect 30168 -6736 30188 -6728
rect 30196 -6736 30224 -6728
rect 30232 -6736 30252 -6728
rect 30288 -6728 30372 -6708
rect 30288 -6736 30308 -6728
rect 30316 -6736 30344 -6728
rect 30352 -6736 30372 -6728
rect 30408 -6728 30492 -6708
rect 30408 -6736 30428 -6728
rect 30436 -6736 30464 -6728
rect 30472 -6736 30492 -6728
rect 30528 -6728 30612 -6708
rect 30528 -6736 30548 -6728
rect 30556 -6736 30584 -6728
rect 30592 -6736 30612 -6728
rect 30648 -6728 30732 -6708
rect 30648 -6736 30668 -6728
rect 30676 -6736 30704 -6728
rect 30712 -6736 30732 -6728
rect 30768 -6728 30852 -6708
rect 30768 -6736 30788 -6728
rect 30796 -6736 30824 -6728
rect 30832 -6736 30852 -6728
rect 30888 -6728 30972 -6708
rect 30888 -6736 30908 -6728
rect 30916 -6736 30944 -6728
rect 30952 -6736 30972 -6728
rect 31008 -6728 31092 -6708
rect 31008 -6736 31028 -6728
rect 31036 -6736 31064 -6728
rect 31072 -6736 31092 -6728
rect 31128 -6728 31212 -6708
rect 31128 -6736 31148 -6728
rect 31156 -6736 31184 -6728
rect 31192 -6736 31212 -6728
rect 31248 -6728 31332 -6708
rect 31248 -6736 31268 -6728
rect 31276 -6736 31304 -6728
rect 31312 -6736 31332 -6728
rect 31368 -6728 31452 -6708
rect 31368 -6736 31388 -6728
rect 31396 -6736 31424 -6728
rect 31432 -6736 31452 -6728
rect 31488 -6728 31572 -6708
rect 31488 -6736 31508 -6728
rect 31516 -6736 31544 -6728
rect 31552 -6736 31572 -6728
rect 31608 -6728 31692 -6708
rect 31608 -6736 31628 -6728
rect 31636 -6736 31664 -6728
rect 31672 -6736 31692 -6728
rect 31728 -6728 31812 -6708
rect 31728 -6736 31748 -6728
rect 31756 -6736 31784 -6728
rect 31792 -6736 31812 -6728
rect 31848 -6728 31932 -6708
rect 31848 -6736 31868 -6728
rect 31876 -6736 31904 -6728
rect 31912 -6736 31932 -6728
rect 31968 -6728 32052 -6708
rect 31968 -6736 31988 -6728
rect 31996 -6736 32024 -6728
rect 32032 -6736 32052 -6728
rect 32088 -6728 32172 -6708
rect 32088 -6736 32108 -6728
rect 32116 -6736 32144 -6728
rect 32152 -6736 32172 -6728
rect 32208 -6728 32292 -6708
rect 32208 -6736 32228 -6728
rect 32236 -6736 32264 -6728
rect 32272 -6736 32292 -6728
rect 32328 -6728 32412 -6708
rect 32328 -6736 32348 -6728
rect 32356 -6736 32384 -6728
rect 32392 -6736 32412 -6728
rect 32448 -6728 32532 -6708
rect 32448 -6736 32468 -6728
rect 32476 -6736 32504 -6728
rect 32512 -6736 32532 -6728
rect 32568 -6728 32652 -6708
rect 32568 -6736 32588 -6728
rect 32596 -6736 32624 -6728
rect 32632 -6736 32652 -6728
rect 32688 -6728 32772 -6708
rect 32688 -6736 32708 -6728
rect 32716 -6736 32744 -6728
rect 32752 -6736 32772 -6728
rect 32808 -6728 32892 -6708
rect 32808 -6736 32828 -6728
rect 32836 -6736 32864 -6728
rect 32872 -6736 32892 -6728
rect 32928 -6728 33012 -6708
rect 32928 -6736 32948 -6728
rect 32956 -6736 32984 -6728
rect 32992 -6736 33012 -6728
rect 33048 -6728 33132 -6708
rect 33048 -6736 33068 -6728
rect 33076 -6736 33104 -6728
rect 33112 -6736 33132 -6728
rect 33168 -6728 33252 -6708
rect 33168 -6736 33188 -6728
rect 33196 -6736 33224 -6728
rect 33232 -6736 33252 -6728
rect 33288 -6728 33372 -6708
rect 33288 -6736 33308 -6728
rect 33316 -6736 33344 -6728
rect 33352 -6736 33372 -6728
rect 33408 -6728 33492 -6708
rect 33408 -6736 33428 -6728
rect 33436 -6736 33464 -6728
rect 33472 -6736 33492 -6728
rect 33528 -6728 33612 -6708
rect 33528 -6736 33548 -6728
rect 33556 -6736 33584 -6728
rect 33592 -6736 33612 -6728
rect 33648 -6728 33732 -6708
rect 33648 -6736 33668 -6728
rect 33676 -6736 33704 -6728
rect 33712 -6736 33732 -6728
rect 33768 -6728 33852 -6708
rect 33768 -6736 33788 -6728
rect 33796 -6736 33824 -6728
rect 33832 -6736 33852 -6728
rect 33888 -6728 33972 -6708
rect 33888 -6736 33908 -6728
rect 33916 -6736 33944 -6728
rect 33952 -6736 33972 -6728
rect 34008 -6728 34092 -6708
rect 34008 -6736 34028 -6728
rect 34036 -6736 34064 -6728
rect 34072 -6736 34092 -6728
rect 34128 -6728 34212 -6708
rect 34128 -6736 34148 -6728
rect 34156 -6736 34184 -6728
rect 34192 -6736 34212 -6728
rect 34248 -6728 34332 -6708
rect 34248 -6736 34268 -6728
rect 34276 -6736 34304 -6728
rect 34312 -6736 34332 -6728
rect 34368 -6728 34452 -6708
rect 34368 -6736 34388 -6728
rect 34396 -6736 34424 -6728
rect 34432 -6736 34452 -6728
rect 34488 -6728 34572 -6708
rect 34488 -6736 34508 -6728
rect 34516 -6736 34544 -6728
rect 34552 -6736 34572 -6728
rect 34608 -6728 34692 -6708
rect 34608 -6736 34628 -6728
rect 34636 -6736 34664 -6728
rect 34672 -6736 34692 -6728
rect 34728 -6728 34812 -6708
rect 34728 -6736 34748 -6728
rect 34756 -6736 34784 -6728
rect 34792 -6736 34812 -6728
rect 34848 -6728 34932 -6708
rect 34848 -6736 34868 -6728
rect 34876 -6736 34904 -6728
rect 34912 -6736 34932 -6728
rect 34968 -6728 35052 -6708
rect 34968 -6736 34988 -6728
rect 34996 -6736 35024 -6728
rect 35032 -6736 35052 -6728
rect 35088 -6728 35172 -6708
rect 35088 -6736 35108 -6728
rect 35116 -6736 35144 -6728
rect 35152 -6736 35172 -6728
rect 35208 -6728 35292 -6708
rect 35208 -6736 35228 -6728
rect 35236 -6736 35264 -6728
rect 35272 -6736 35292 -6728
rect 35328 -6728 35412 -6708
rect 35328 -6736 35348 -6728
rect 35356 -6736 35384 -6728
rect 35392 -6736 35412 -6728
rect 35448 -6728 35532 -6708
rect 35448 -6736 35468 -6728
rect 35476 -6736 35504 -6728
rect 35512 -6736 35532 -6728
rect 35568 -6728 35652 -6708
rect 35568 -6736 35588 -6728
rect 35596 -6736 35624 -6728
rect 35632 -6736 35652 -6728
rect 35688 -6728 35772 -6708
rect 35688 -6736 35708 -6728
rect 35716 -6736 35744 -6728
rect 35752 -6736 35772 -6728
rect 35808 -6728 35892 -6708
rect 35808 -6736 35828 -6728
rect 35836 -6736 35864 -6728
rect 35872 -6736 35892 -6728
rect 35928 -6728 36012 -6708
rect 35928 -6736 35948 -6728
rect 35956 -6736 35984 -6728
rect 35992 -6736 36012 -6728
rect 36048 -6728 36132 -6708
rect 36048 -6736 36068 -6728
rect 36076 -6736 36104 -6728
rect 36112 -6736 36132 -6728
rect 36168 -6728 36252 -6708
rect 36168 -6736 36188 -6728
rect 36196 -6736 36224 -6728
rect 36232 -6736 36252 -6728
rect 36288 -6728 36372 -6708
rect 36288 -6736 36308 -6728
rect 36316 -6736 36344 -6728
rect 36352 -6736 36372 -6728
rect 36408 -6728 36492 -6708
rect 36408 -6736 36428 -6728
rect 36436 -6736 36464 -6728
rect 36472 -6736 36492 -6728
rect 36528 -6728 36612 -6708
rect 36528 -6736 36548 -6728
rect 36556 -6736 36584 -6728
rect 36592 -6736 36612 -6728
rect 36648 -6728 36732 -6708
rect 36648 -6736 36668 -6728
rect 36676 -6736 36704 -6728
rect 36712 -6736 36732 -6728
rect 36768 -6728 36852 -6708
rect 36768 -6736 36788 -6728
rect 36796 -6736 36824 -6728
rect 36832 -6736 36852 -6728
rect 36888 -6728 36972 -6708
rect 36888 -6736 36908 -6728
rect 36916 -6736 36944 -6728
rect 36952 -6736 36972 -6728
rect 37008 -6728 37092 -6708
rect 37008 -6736 37028 -6728
rect 37036 -6736 37064 -6728
rect 37072 -6736 37092 -6728
rect 37128 -6728 37212 -6708
rect 37128 -6736 37148 -6728
rect 37156 -6736 37184 -6728
rect 37192 -6736 37212 -6728
rect 37248 -6728 37332 -6708
rect 37248 -6736 37268 -6728
rect 37276 -6736 37304 -6728
rect 37312 -6736 37332 -6728
rect 37368 -6728 37452 -6708
rect 37368 -6736 37388 -6728
rect 37396 -6736 37424 -6728
rect 37432 -6736 37452 -6728
rect 37488 -6728 37572 -6708
rect 37488 -6736 37508 -6728
rect 37516 -6736 37544 -6728
rect 37552 -6736 37572 -6728
rect 37608 -6728 37692 -6708
rect 37608 -6736 37628 -6728
rect 37636 -6736 37664 -6728
rect 37672 -6736 37692 -6728
rect 37728 -6728 37812 -6708
rect 37728 -6736 37748 -6728
rect 37756 -6736 37784 -6728
rect 37792 -6736 37812 -6728
rect 37848 -6728 37932 -6708
rect 37848 -6736 37868 -6728
rect 37876 -6736 37904 -6728
rect 37912 -6736 37932 -6728
rect 37968 -6728 38052 -6708
rect 37968 -6736 37988 -6728
rect 37996 -6736 38024 -6728
rect 38032 -6736 38052 -6728
rect 38088 -6728 38172 -6708
rect 38088 -6736 38108 -6728
rect 38116 -6736 38144 -6728
rect 38152 -6736 38172 -6728
rect 38208 -6728 38292 -6708
rect 38208 -6736 38228 -6728
rect 38236 -6736 38264 -6728
rect 38272 -6736 38292 -6728
rect 38328 -6728 38412 -6708
rect 38328 -6736 38348 -6728
rect 38356 -6736 38384 -6728
rect 38392 -6736 38412 -6728
rect 38448 -6728 38532 -6708
rect 38448 -6736 38468 -6728
rect 38476 -6736 38504 -6728
rect 38512 -6736 38532 -6728
rect 38568 -6728 38652 -6708
rect 38568 -6736 38588 -6728
rect 38596 -6736 38624 -6728
rect 38632 -6736 38652 -6728
rect 38688 -6728 38772 -6708
rect 38688 -6736 38708 -6728
rect 38716 -6736 38744 -6728
rect 38752 -6736 38772 -6728
rect 38808 -6728 38892 -6708
rect 38808 -6736 38828 -6728
rect 38836 -6736 38864 -6728
rect 38872 -6736 38892 -6728
rect 38928 -6728 39012 -6708
rect 38928 -6736 38948 -6728
rect 38956 -6736 38984 -6728
rect 38992 -6736 39012 -6728
rect 39048 -6728 39132 -6708
rect 39048 -6736 39068 -6728
rect 39076 -6736 39104 -6728
rect 39112 -6736 39132 -6728
rect 39168 -6728 39252 -6708
rect 39168 -6736 39188 -6728
rect 39196 -6736 39224 -6728
rect 39232 -6736 39252 -6728
rect 39288 -6728 39372 -6708
rect 39288 -6736 39308 -6728
rect 39316 -6736 39344 -6728
rect 39352 -6736 39372 -6728
rect 39408 -6728 39492 -6708
rect 39408 -6736 39428 -6728
rect 39436 -6736 39464 -6728
rect 39472 -6736 39492 -6728
rect 39528 -6728 39612 -6708
rect 39528 -6736 39548 -6728
rect 39556 -6736 39584 -6728
rect 39592 -6736 39612 -6728
rect 39648 -6728 39732 -6708
rect 39648 -6736 39668 -6728
rect 39676 -6736 39704 -6728
rect 39712 -6736 39732 -6728
rect 39768 -6728 39852 -6708
rect 39768 -6736 39788 -6728
rect 39796 -6736 39824 -6728
rect 39832 -6736 39852 -6728
rect 39888 -6728 39972 -6708
rect 39888 -6736 39908 -6728
rect 39916 -6736 39944 -6728
rect 39952 -6736 39972 -6728
rect 40008 -6728 40092 -6708
rect 40008 -6736 40028 -6728
rect 40036 -6736 40064 -6728
rect 40072 -6736 40092 -6728
rect 40128 -6728 40212 -6708
rect 40128 -6736 40148 -6728
rect 40156 -6736 40184 -6728
rect 40192 -6736 40212 -6728
rect 40248 -6728 40332 -6708
rect 40248 -6736 40268 -6728
rect 40276 -6736 40304 -6728
rect 40312 -6736 40332 -6728
rect 40368 -6728 40452 -6708
rect 40368 -6736 40388 -6728
rect 40396 -6736 40424 -6728
rect 40432 -6736 40452 -6728
rect 40488 -6728 40572 -6708
rect 40488 -6736 40508 -6728
rect 40516 -6736 40544 -6728
rect 40552 -6736 40572 -6728
rect 40608 -6728 40692 -6708
rect 40608 -6736 40628 -6728
rect 40636 -6736 40664 -6728
rect 40672 -6736 40692 -6728
rect 40728 -6728 40812 -6708
rect 40728 -6736 40748 -6728
rect 40756 -6736 40784 -6728
rect 40792 -6736 40812 -6728
rect 40848 -6728 40932 -6708
rect 40848 -6736 40868 -6728
rect 40876 -6736 40904 -6728
rect 40912 -6736 40932 -6728
rect 40968 -6728 41052 -6708
rect 40968 -6736 40988 -6728
rect 40996 -6736 41024 -6728
rect 41032 -6736 41052 -6728
rect 41088 -6728 41172 -6708
rect 41088 -6736 41108 -6728
rect 41116 -6736 41144 -6728
rect 41152 -6736 41172 -6728
rect 41208 -6728 41292 -6708
rect 41208 -6736 41228 -6728
rect 41236 -6736 41264 -6728
rect 41272 -6736 41292 -6728
rect 41328 -6728 41412 -6708
rect 41328 -6736 41348 -6728
rect 41356 -6736 41384 -6728
rect 41392 -6736 41412 -6728
rect 41448 -6728 41532 -6708
rect 41448 -6736 41468 -6728
rect 41476 -6736 41504 -6728
rect 41512 -6736 41532 -6728
rect 41568 -6728 41652 -6708
rect 41568 -6736 41588 -6728
rect 41596 -6736 41624 -6728
rect 41632 -6736 41652 -6728
rect 41688 -6728 41772 -6708
rect 41688 -6736 41708 -6728
rect 41716 -6736 41744 -6728
rect 41752 -6736 41772 -6728
rect 41808 -6728 41892 -6708
rect 41808 -6736 41828 -6728
rect 41836 -6736 41864 -6728
rect 41872 -6736 41892 -6728
rect 41928 -6728 42012 -6708
rect 41928 -6736 41948 -6728
rect 41956 -6736 41984 -6728
rect 41992 -6736 42012 -6728
rect 42048 -6728 42132 -6708
rect 42048 -6736 42068 -6728
rect 42076 -6736 42104 -6728
rect 42112 -6736 42132 -6728
rect 42168 -6728 42252 -6708
rect 42168 -6736 42188 -6728
rect 42196 -6736 42224 -6728
rect 42232 -6736 42252 -6728
rect 42288 -6728 42372 -6708
rect 42288 -6736 42308 -6728
rect 42316 -6736 42344 -6728
rect 42352 -6736 42372 -6728
rect 42408 -6728 42492 -6708
rect 42408 -6736 42428 -6728
rect 42436 -6736 42464 -6728
rect 42472 -6736 42492 -6728
rect 42528 -6728 42612 -6708
rect 42528 -6736 42548 -6728
rect 42556 -6736 42584 -6728
rect 42592 -6736 42612 -6728
rect 42648 -6728 42732 -6708
rect 42648 -6736 42668 -6728
rect 42676 -6736 42704 -6728
rect 42712 -6736 42732 -6728
rect 42768 -6728 42852 -6708
rect 42768 -6736 42788 -6728
rect 42796 -6736 42824 -6728
rect 42832 -6736 42852 -6728
rect 42888 -6728 42972 -6708
rect 42888 -6736 42908 -6728
rect 42916 -6736 42944 -6728
rect 42952 -6736 42972 -6728
rect 43008 -6728 43092 -6708
rect 43008 -6736 43028 -6728
rect 43036 -6736 43064 -6728
rect 43072 -6736 43092 -6728
rect 43128 -6728 43212 -6708
rect 43128 -6736 43148 -6728
rect 43156 -6736 43184 -6728
rect 43192 -6736 43212 -6728
rect 43248 -6728 43332 -6708
rect 43248 -6736 43268 -6728
rect 43276 -6736 43304 -6728
rect 43312 -6736 43332 -6728
rect 43368 -6728 43452 -6708
rect 43368 -6736 43388 -6728
rect 43396 -6736 43424 -6728
rect 43432 -6736 43452 -6728
rect 43488 -6728 43572 -6708
rect 43488 -6736 43508 -6728
rect 43516 -6736 43544 -6728
rect 43552 -6736 43572 -6728
rect 43608 -6728 43692 -6708
rect 43608 -6736 43628 -6728
rect 43636 -6736 43664 -6728
rect 43672 -6736 43692 -6728
rect 43728 -6728 43812 -6708
rect 43728 -6736 43748 -6728
rect 43756 -6736 43784 -6728
rect 43792 -6736 43812 -6728
rect 43848 -6728 43932 -6708
rect 43848 -6736 43868 -6728
rect 43876 -6736 43904 -6728
rect 43912 -6736 43932 -6728
rect 43968 -6728 44052 -6708
rect 43968 -6736 43988 -6728
rect 43996 -6736 44024 -6728
rect 44032 -6736 44052 -6728
rect 44088 -6728 44172 -6708
rect 44088 -6736 44108 -6728
rect 44116 -6736 44144 -6728
rect 44152 -6736 44172 -6728
rect 44208 -6728 44292 -6708
rect 44208 -6736 44228 -6728
rect 44236 -6736 44264 -6728
rect 44272 -6736 44292 -6728
rect 44328 -6728 44412 -6708
rect 44328 -6736 44348 -6728
rect 44356 -6736 44384 -6728
rect 44392 -6736 44412 -6728
rect 44448 -6728 44532 -6708
rect 44448 -6736 44468 -6728
rect 44476 -6736 44504 -6728
rect 44512 -6736 44532 -6728
rect 44568 -6728 44652 -6708
rect 44568 -6736 44588 -6728
rect 44596 -6736 44624 -6728
rect 44632 -6736 44652 -6728
rect 44688 -6728 44772 -6708
rect 44688 -6736 44708 -6728
rect 44716 -6736 44744 -6728
rect 44752 -6736 44772 -6728
rect 44808 -6728 44892 -6708
rect 44808 -6736 44828 -6728
rect 44836 -6736 44864 -6728
rect 44872 -6736 44892 -6728
rect 44928 -6728 45012 -6708
rect 44928 -6736 44948 -6728
rect 44956 -6736 44984 -6728
rect 44992 -6736 45012 -6728
rect 45048 -6728 45132 -6708
rect 45048 -6736 45068 -6728
rect 45076 -6736 45104 -6728
rect 45112 -6736 45132 -6728
rect 45168 -6728 45252 -6708
rect 45168 -6736 45188 -6728
rect 45196 -6736 45224 -6728
rect 45232 -6736 45252 -6728
rect 45288 -6728 45372 -6708
rect 45288 -6736 45308 -6728
rect 45316 -6736 45344 -6728
rect 45352 -6736 45372 -6728
rect 45408 -6728 45492 -6708
rect 45408 -6736 45428 -6728
rect 45436 -6736 45464 -6728
rect 45472 -6736 45492 -6728
rect 45528 -6728 45612 -6708
rect 45528 -6736 45548 -6728
rect 45556 -6736 45584 -6728
rect 45592 -6736 45612 -6728
rect 25876 -6764 25932 -6736
rect 25996 -6764 26052 -6736
rect 26116 -6764 26172 -6736
rect 26236 -6764 26292 -6736
rect 26356 -6764 26412 -6736
rect 26476 -6764 26532 -6736
rect 26596 -6764 26652 -6736
rect 26716 -6764 26772 -6736
rect 26836 -6764 26892 -6736
rect 26956 -6764 27012 -6736
rect 27076 -6764 27132 -6736
rect 27196 -6764 27252 -6736
rect 27316 -6764 27372 -6736
rect 27436 -6764 27492 -6736
rect 27556 -6764 27612 -6736
rect 27676 -6764 27732 -6736
rect 27796 -6764 27852 -6736
rect 27916 -6764 27972 -6736
rect 28036 -6764 28092 -6736
rect 28156 -6764 28212 -6736
rect 28276 -6764 28332 -6736
rect 28396 -6764 28452 -6736
rect 28516 -6764 28572 -6736
rect 28636 -6764 28692 -6736
rect 28756 -6764 28812 -6736
rect 28876 -6764 28932 -6736
rect 28996 -6764 29052 -6736
rect 29116 -6764 29172 -6736
rect 29236 -6764 29292 -6736
rect 29356 -6764 29412 -6736
rect 29476 -6764 29532 -6736
rect 29596 -6764 29652 -6736
rect 29716 -6764 29772 -6736
rect 29836 -6764 29892 -6736
rect 29956 -6764 30012 -6736
rect 30076 -6764 30132 -6736
rect 30196 -6764 30252 -6736
rect 30316 -6764 30372 -6736
rect 30436 -6764 30492 -6736
rect 30556 -6764 30612 -6736
rect 30676 -6764 30732 -6736
rect 30796 -6764 30852 -6736
rect 30916 -6764 30972 -6736
rect 31036 -6764 31092 -6736
rect 31156 -6764 31212 -6736
rect 31276 -6764 31332 -6736
rect 31396 -6764 31452 -6736
rect 31516 -6764 31572 -6736
rect 31636 -6764 31692 -6736
rect 31756 -6764 31812 -6736
rect 31876 -6764 31932 -6736
rect 31996 -6764 32052 -6736
rect 32116 -6764 32172 -6736
rect 32236 -6764 32292 -6736
rect 32356 -6764 32412 -6736
rect 32476 -6764 32532 -6736
rect 32596 -6764 32652 -6736
rect 32716 -6764 32772 -6736
rect 32836 -6764 32892 -6736
rect 32956 -6764 33012 -6736
rect 33076 -6764 33132 -6736
rect 33196 -6764 33252 -6736
rect 33316 -6764 33372 -6736
rect 33436 -6764 33492 -6736
rect 33556 -6764 33612 -6736
rect 33676 -6764 33732 -6736
rect 33796 -6764 33852 -6736
rect 33916 -6764 33972 -6736
rect 34036 -6764 34092 -6736
rect 34156 -6764 34212 -6736
rect 34276 -6764 34332 -6736
rect 34396 -6764 34452 -6736
rect 34516 -6764 34572 -6736
rect 34636 -6764 34692 -6736
rect 34756 -6764 34812 -6736
rect 34876 -6764 34932 -6736
rect 34996 -6764 35052 -6736
rect 35116 -6764 35172 -6736
rect 35236 -6764 35292 -6736
rect 35356 -6764 35412 -6736
rect 35476 -6764 35532 -6736
rect 35596 -6764 35652 -6736
rect 35716 -6764 35772 -6736
rect 35836 -6764 35892 -6736
rect 35956 -6764 36012 -6736
rect 36076 -6764 36132 -6736
rect 36196 -6764 36252 -6736
rect 36316 -6764 36372 -6736
rect 36436 -6764 36492 -6736
rect 36556 -6764 36612 -6736
rect 36676 -6764 36732 -6736
rect 36796 -6764 36852 -6736
rect 36916 -6764 36972 -6736
rect 37036 -6764 37092 -6736
rect 37156 -6764 37212 -6736
rect 37276 -6764 37332 -6736
rect 37396 -6764 37452 -6736
rect 37516 -6764 37572 -6736
rect 37636 -6764 37692 -6736
rect 37756 -6764 37812 -6736
rect 37876 -6764 37932 -6736
rect 37996 -6764 38052 -6736
rect 38116 -6764 38172 -6736
rect 38236 -6764 38292 -6736
rect 38356 -6764 38412 -6736
rect 38476 -6764 38532 -6736
rect 38596 -6764 38652 -6736
rect 38716 -6764 38772 -6736
rect 38836 -6764 38892 -6736
rect 38956 -6764 39012 -6736
rect 39076 -6764 39132 -6736
rect 39196 -6764 39252 -6736
rect 39316 -6764 39372 -6736
rect 39436 -6764 39492 -6736
rect 39556 -6764 39612 -6736
rect 39676 -6764 39732 -6736
rect 39796 -6764 39852 -6736
rect 39916 -6764 39972 -6736
rect 40036 -6764 40092 -6736
rect 40156 -6764 40212 -6736
rect 40276 -6764 40332 -6736
rect 40396 -6764 40452 -6736
rect 40516 -6764 40572 -6736
rect 40636 -6764 40692 -6736
rect 40756 -6764 40812 -6736
rect 40876 -6764 40932 -6736
rect 40996 -6764 41052 -6736
rect 41116 -6764 41172 -6736
rect 41236 -6764 41292 -6736
rect 41356 -6764 41412 -6736
rect 41476 -6764 41532 -6736
rect 41596 -6764 41652 -6736
rect 41716 -6764 41772 -6736
rect 41836 -6764 41892 -6736
rect 41956 -6764 42012 -6736
rect 42076 -6764 42132 -6736
rect 42196 -6764 42252 -6736
rect 42316 -6764 42372 -6736
rect 42436 -6764 42492 -6736
rect 42556 -6764 42612 -6736
rect 42676 -6764 42732 -6736
rect 42796 -6764 42852 -6736
rect 42916 -6764 42972 -6736
rect 43036 -6764 43092 -6736
rect 43156 -6764 43212 -6736
rect 43276 -6764 43332 -6736
rect 43396 -6764 43452 -6736
rect 43516 -6764 43572 -6736
rect 43636 -6764 43692 -6736
rect 43756 -6764 43812 -6736
rect 43876 -6764 43932 -6736
rect 43996 -6764 44052 -6736
rect 44116 -6764 44172 -6736
rect 44236 -6764 44292 -6736
rect 44356 -6764 44412 -6736
rect 44476 -6764 44532 -6736
rect 44596 -6764 44652 -6736
rect 44716 -6764 44772 -6736
rect 44836 -6764 44892 -6736
rect 44956 -6764 45012 -6736
rect 45076 -6764 45132 -6736
rect 45196 -6764 45252 -6736
rect 45316 -6764 45372 -6736
rect 45436 -6764 45492 -6736
rect 45556 -6764 45612 -6736
rect 25848 -6908 25932 -6888
rect 25848 -6916 25868 -6908
rect 25876 -6916 25904 -6908
rect 25912 -6916 25932 -6908
rect 25968 -6908 26052 -6888
rect 25968 -6916 25988 -6908
rect 25996 -6916 26024 -6908
rect 26032 -6916 26052 -6908
rect 26088 -6908 26172 -6888
rect 26088 -6916 26108 -6908
rect 26116 -6916 26144 -6908
rect 26152 -6916 26172 -6908
rect 26208 -6908 26292 -6888
rect 26208 -6916 26228 -6908
rect 26236 -6916 26264 -6908
rect 26272 -6916 26292 -6908
rect 26328 -6908 26412 -6888
rect 26328 -6916 26348 -6908
rect 26356 -6916 26384 -6908
rect 26392 -6916 26412 -6908
rect 26448 -6908 26532 -6888
rect 26448 -6916 26468 -6908
rect 26476 -6916 26504 -6908
rect 26512 -6916 26532 -6908
rect 26568 -6908 26652 -6888
rect 26568 -6916 26588 -6908
rect 26596 -6916 26624 -6908
rect 26632 -6916 26652 -6908
rect 26688 -6908 26772 -6888
rect 26688 -6916 26708 -6908
rect 26716 -6916 26744 -6908
rect 26752 -6916 26772 -6908
rect 26808 -6908 26892 -6888
rect 26808 -6916 26828 -6908
rect 26836 -6916 26864 -6908
rect 26872 -6916 26892 -6908
rect 26928 -6908 27012 -6888
rect 26928 -6916 26948 -6908
rect 26956 -6916 26984 -6908
rect 26992 -6916 27012 -6908
rect 27048 -6908 27132 -6888
rect 27048 -6916 27068 -6908
rect 27076 -6916 27104 -6908
rect 27112 -6916 27132 -6908
rect 27168 -6908 27252 -6888
rect 27168 -6916 27188 -6908
rect 27196 -6916 27224 -6908
rect 27232 -6916 27252 -6908
rect 27288 -6908 27372 -6888
rect 27288 -6916 27308 -6908
rect 27316 -6916 27344 -6908
rect 27352 -6916 27372 -6908
rect 27408 -6908 27492 -6888
rect 27408 -6916 27428 -6908
rect 27436 -6916 27464 -6908
rect 27472 -6916 27492 -6908
rect 27528 -6908 27612 -6888
rect 27528 -6916 27548 -6908
rect 27556 -6916 27584 -6908
rect 27592 -6916 27612 -6908
rect 27648 -6908 27732 -6888
rect 27648 -6916 27668 -6908
rect 27676 -6916 27704 -6908
rect 27712 -6916 27732 -6908
rect 27768 -6908 27852 -6888
rect 27768 -6916 27788 -6908
rect 27796 -6916 27824 -6908
rect 27832 -6916 27852 -6908
rect 27888 -6908 27972 -6888
rect 27888 -6916 27908 -6908
rect 27916 -6916 27944 -6908
rect 27952 -6916 27972 -6908
rect 28008 -6908 28092 -6888
rect 28008 -6916 28028 -6908
rect 28036 -6916 28064 -6908
rect 28072 -6916 28092 -6908
rect 28128 -6908 28212 -6888
rect 28128 -6916 28148 -6908
rect 28156 -6916 28184 -6908
rect 28192 -6916 28212 -6908
rect 28248 -6908 28332 -6888
rect 28248 -6916 28268 -6908
rect 28276 -6916 28304 -6908
rect 28312 -6916 28332 -6908
rect 28368 -6908 28452 -6888
rect 28368 -6916 28388 -6908
rect 28396 -6916 28424 -6908
rect 28432 -6916 28452 -6908
rect 28488 -6908 28572 -6888
rect 28488 -6916 28508 -6908
rect 28516 -6916 28544 -6908
rect 28552 -6916 28572 -6908
rect 28608 -6908 28692 -6888
rect 28608 -6916 28628 -6908
rect 28636 -6916 28664 -6908
rect 28672 -6916 28692 -6908
rect 28728 -6908 28812 -6888
rect 28728 -6916 28748 -6908
rect 28756 -6916 28784 -6908
rect 28792 -6916 28812 -6908
rect 28848 -6908 28932 -6888
rect 28848 -6916 28868 -6908
rect 28876 -6916 28904 -6908
rect 28912 -6916 28932 -6908
rect 28968 -6908 29052 -6888
rect 28968 -6916 28988 -6908
rect 28996 -6916 29024 -6908
rect 29032 -6916 29052 -6908
rect 29088 -6908 29172 -6888
rect 29088 -6916 29108 -6908
rect 29116 -6916 29144 -6908
rect 29152 -6916 29172 -6908
rect 29208 -6908 29292 -6888
rect 29208 -6916 29228 -6908
rect 29236 -6916 29264 -6908
rect 29272 -6916 29292 -6908
rect 29328 -6908 29412 -6888
rect 29328 -6916 29348 -6908
rect 29356 -6916 29384 -6908
rect 29392 -6916 29412 -6908
rect 29448 -6908 29532 -6888
rect 29448 -6916 29468 -6908
rect 29476 -6916 29504 -6908
rect 29512 -6916 29532 -6908
rect 29568 -6908 29652 -6888
rect 29568 -6916 29588 -6908
rect 29596 -6916 29624 -6908
rect 29632 -6916 29652 -6908
rect 29688 -6908 29772 -6888
rect 29688 -6916 29708 -6908
rect 29716 -6916 29744 -6908
rect 29752 -6916 29772 -6908
rect 29808 -6908 29892 -6888
rect 29808 -6916 29828 -6908
rect 29836 -6916 29864 -6908
rect 29872 -6916 29892 -6908
rect 29928 -6908 30012 -6888
rect 29928 -6916 29948 -6908
rect 29956 -6916 29984 -6908
rect 29992 -6916 30012 -6908
rect 30048 -6908 30132 -6888
rect 30048 -6916 30068 -6908
rect 30076 -6916 30104 -6908
rect 30112 -6916 30132 -6908
rect 30168 -6908 30252 -6888
rect 30168 -6916 30188 -6908
rect 30196 -6916 30224 -6908
rect 30232 -6916 30252 -6908
rect 30288 -6908 30372 -6888
rect 30288 -6916 30308 -6908
rect 30316 -6916 30344 -6908
rect 30352 -6916 30372 -6908
rect 30408 -6908 30492 -6888
rect 30408 -6916 30428 -6908
rect 30436 -6916 30464 -6908
rect 30472 -6916 30492 -6908
rect 30528 -6908 30612 -6888
rect 30528 -6916 30548 -6908
rect 30556 -6916 30584 -6908
rect 30592 -6916 30612 -6908
rect 30648 -6908 30732 -6888
rect 30648 -6916 30668 -6908
rect 30676 -6916 30704 -6908
rect 30712 -6916 30732 -6908
rect 30768 -6908 30852 -6888
rect 30768 -6916 30788 -6908
rect 30796 -6916 30824 -6908
rect 30832 -6916 30852 -6908
rect 30888 -6908 30972 -6888
rect 30888 -6916 30908 -6908
rect 30916 -6916 30944 -6908
rect 30952 -6916 30972 -6908
rect 31008 -6908 31092 -6888
rect 31008 -6916 31028 -6908
rect 31036 -6916 31064 -6908
rect 31072 -6916 31092 -6908
rect 31128 -6908 31212 -6888
rect 31128 -6916 31148 -6908
rect 31156 -6916 31184 -6908
rect 31192 -6916 31212 -6908
rect 31248 -6908 31332 -6888
rect 31248 -6916 31268 -6908
rect 31276 -6916 31304 -6908
rect 31312 -6916 31332 -6908
rect 31368 -6908 31452 -6888
rect 31368 -6916 31388 -6908
rect 31396 -6916 31424 -6908
rect 31432 -6916 31452 -6908
rect 31488 -6908 31572 -6888
rect 31488 -6916 31508 -6908
rect 31516 -6916 31544 -6908
rect 31552 -6916 31572 -6908
rect 31608 -6908 31692 -6888
rect 31608 -6916 31628 -6908
rect 31636 -6916 31664 -6908
rect 31672 -6916 31692 -6908
rect 31728 -6908 31812 -6888
rect 31728 -6916 31748 -6908
rect 31756 -6916 31784 -6908
rect 31792 -6916 31812 -6908
rect 31848 -6908 31932 -6888
rect 31848 -6916 31868 -6908
rect 31876 -6916 31904 -6908
rect 31912 -6916 31932 -6908
rect 31968 -6908 32052 -6888
rect 31968 -6916 31988 -6908
rect 31996 -6916 32024 -6908
rect 32032 -6916 32052 -6908
rect 32088 -6908 32172 -6888
rect 32088 -6916 32108 -6908
rect 32116 -6916 32144 -6908
rect 32152 -6916 32172 -6908
rect 32208 -6908 32292 -6888
rect 32208 -6916 32228 -6908
rect 32236 -6916 32264 -6908
rect 32272 -6916 32292 -6908
rect 32328 -6908 32412 -6888
rect 32328 -6916 32348 -6908
rect 32356 -6916 32384 -6908
rect 32392 -6916 32412 -6908
rect 32448 -6908 32532 -6888
rect 32448 -6916 32468 -6908
rect 32476 -6916 32504 -6908
rect 32512 -6916 32532 -6908
rect 32568 -6908 32652 -6888
rect 32568 -6916 32588 -6908
rect 32596 -6916 32624 -6908
rect 32632 -6916 32652 -6908
rect 32688 -6908 32772 -6888
rect 32688 -6916 32708 -6908
rect 32716 -6916 32744 -6908
rect 32752 -6916 32772 -6908
rect 32808 -6908 32892 -6888
rect 32808 -6916 32828 -6908
rect 32836 -6916 32864 -6908
rect 32872 -6916 32892 -6908
rect 32928 -6908 33012 -6888
rect 32928 -6916 32948 -6908
rect 32956 -6916 32984 -6908
rect 32992 -6916 33012 -6908
rect 33048 -6908 33132 -6888
rect 33048 -6916 33068 -6908
rect 33076 -6916 33104 -6908
rect 33112 -6916 33132 -6908
rect 33168 -6908 33252 -6888
rect 33168 -6916 33188 -6908
rect 33196 -6916 33224 -6908
rect 33232 -6916 33252 -6908
rect 33288 -6908 33372 -6888
rect 33288 -6916 33308 -6908
rect 33316 -6916 33344 -6908
rect 33352 -6916 33372 -6908
rect 33408 -6908 33492 -6888
rect 33408 -6916 33428 -6908
rect 33436 -6916 33464 -6908
rect 33472 -6916 33492 -6908
rect 33528 -6908 33612 -6888
rect 33528 -6916 33548 -6908
rect 33556 -6916 33584 -6908
rect 33592 -6916 33612 -6908
rect 33648 -6908 33732 -6888
rect 33648 -6916 33668 -6908
rect 33676 -6916 33704 -6908
rect 33712 -6916 33732 -6908
rect 33768 -6908 33852 -6888
rect 33768 -6916 33788 -6908
rect 33796 -6916 33824 -6908
rect 33832 -6916 33852 -6908
rect 33888 -6908 33972 -6888
rect 33888 -6916 33908 -6908
rect 33916 -6916 33944 -6908
rect 33952 -6916 33972 -6908
rect 34008 -6908 34092 -6888
rect 34008 -6916 34028 -6908
rect 34036 -6916 34064 -6908
rect 34072 -6916 34092 -6908
rect 34128 -6908 34212 -6888
rect 34128 -6916 34148 -6908
rect 34156 -6916 34184 -6908
rect 34192 -6916 34212 -6908
rect 34248 -6908 34332 -6888
rect 34248 -6916 34268 -6908
rect 34276 -6916 34304 -6908
rect 34312 -6916 34332 -6908
rect 34368 -6908 34452 -6888
rect 34368 -6916 34388 -6908
rect 34396 -6916 34424 -6908
rect 34432 -6916 34452 -6908
rect 34488 -6908 34572 -6888
rect 34488 -6916 34508 -6908
rect 34516 -6916 34544 -6908
rect 34552 -6916 34572 -6908
rect 34608 -6908 34692 -6888
rect 34608 -6916 34628 -6908
rect 34636 -6916 34664 -6908
rect 34672 -6916 34692 -6908
rect 34728 -6908 34812 -6888
rect 34728 -6916 34748 -6908
rect 34756 -6916 34784 -6908
rect 34792 -6916 34812 -6908
rect 34848 -6908 34932 -6888
rect 34848 -6916 34868 -6908
rect 34876 -6916 34904 -6908
rect 34912 -6916 34932 -6908
rect 34968 -6908 35052 -6888
rect 34968 -6916 34988 -6908
rect 34996 -6916 35024 -6908
rect 35032 -6916 35052 -6908
rect 35088 -6908 35172 -6888
rect 35088 -6916 35108 -6908
rect 35116 -6916 35144 -6908
rect 35152 -6916 35172 -6908
rect 35208 -6908 35292 -6888
rect 35208 -6916 35228 -6908
rect 35236 -6916 35264 -6908
rect 35272 -6916 35292 -6908
rect 35328 -6908 35412 -6888
rect 35328 -6916 35348 -6908
rect 35356 -6916 35384 -6908
rect 35392 -6916 35412 -6908
rect 35448 -6908 35532 -6888
rect 35448 -6916 35468 -6908
rect 35476 -6916 35504 -6908
rect 35512 -6916 35532 -6908
rect 35568 -6908 35652 -6888
rect 35568 -6916 35588 -6908
rect 35596 -6916 35624 -6908
rect 35632 -6916 35652 -6908
rect 35688 -6908 35772 -6888
rect 35688 -6916 35708 -6908
rect 35716 -6916 35744 -6908
rect 35752 -6916 35772 -6908
rect 35808 -6908 35892 -6888
rect 35808 -6916 35828 -6908
rect 35836 -6916 35864 -6908
rect 35872 -6916 35892 -6908
rect 35928 -6908 36012 -6888
rect 35928 -6916 35948 -6908
rect 35956 -6916 35984 -6908
rect 35992 -6916 36012 -6908
rect 36048 -6908 36132 -6888
rect 36048 -6916 36068 -6908
rect 36076 -6916 36104 -6908
rect 36112 -6916 36132 -6908
rect 36168 -6908 36252 -6888
rect 36168 -6916 36188 -6908
rect 36196 -6916 36224 -6908
rect 36232 -6916 36252 -6908
rect 36288 -6908 36372 -6888
rect 36288 -6916 36308 -6908
rect 36316 -6916 36344 -6908
rect 36352 -6916 36372 -6908
rect 36408 -6908 36492 -6888
rect 36408 -6916 36428 -6908
rect 36436 -6916 36464 -6908
rect 36472 -6916 36492 -6908
rect 36528 -6908 36612 -6888
rect 36528 -6916 36548 -6908
rect 36556 -6916 36584 -6908
rect 36592 -6916 36612 -6908
rect 36648 -6908 36732 -6888
rect 36648 -6916 36668 -6908
rect 36676 -6916 36704 -6908
rect 36712 -6916 36732 -6908
rect 36768 -6908 36852 -6888
rect 36768 -6916 36788 -6908
rect 36796 -6916 36824 -6908
rect 36832 -6916 36852 -6908
rect 36888 -6908 36972 -6888
rect 36888 -6916 36908 -6908
rect 36916 -6916 36944 -6908
rect 36952 -6916 36972 -6908
rect 37008 -6908 37092 -6888
rect 37008 -6916 37028 -6908
rect 37036 -6916 37064 -6908
rect 37072 -6916 37092 -6908
rect 37128 -6908 37212 -6888
rect 37128 -6916 37148 -6908
rect 37156 -6916 37184 -6908
rect 37192 -6916 37212 -6908
rect 37248 -6908 37332 -6888
rect 37248 -6916 37268 -6908
rect 37276 -6916 37304 -6908
rect 37312 -6916 37332 -6908
rect 37368 -6908 37452 -6888
rect 37368 -6916 37388 -6908
rect 37396 -6916 37424 -6908
rect 37432 -6916 37452 -6908
rect 37488 -6908 37572 -6888
rect 37488 -6916 37508 -6908
rect 37516 -6916 37544 -6908
rect 37552 -6916 37572 -6908
rect 37608 -6908 37692 -6888
rect 37608 -6916 37628 -6908
rect 37636 -6916 37664 -6908
rect 37672 -6916 37692 -6908
rect 37728 -6908 37812 -6888
rect 37728 -6916 37748 -6908
rect 37756 -6916 37784 -6908
rect 37792 -6916 37812 -6908
rect 37848 -6908 37932 -6888
rect 37848 -6916 37868 -6908
rect 37876 -6916 37904 -6908
rect 37912 -6916 37932 -6908
rect 37968 -6908 38052 -6888
rect 37968 -6916 37988 -6908
rect 37996 -6916 38024 -6908
rect 38032 -6916 38052 -6908
rect 38088 -6908 38172 -6888
rect 38088 -6916 38108 -6908
rect 38116 -6916 38144 -6908
rect 38152 -6916 38172 -6908
rect 38208 -6908 38292 -6888
rect 38208 -6916 38228 -6908
rect 38236 -6916 38264 -6908
rect 38272 -6916 38292 -6908
rect 38328 -6908 38412 -6888
rect 38328 -6916 38348 -6908
rect 38356 -6916 38384 -6908
rect 38392 -6916 38412 -6908
rect 38448 -6908 38532 -6888
rect 38448 -6916 38468 -6908
rect 38476 -6916 38504 -6908
rect 38512 -6916 38532 -6908
rect 38568 -6908 38652 -6888
rect 38568 -6916 38588 -6908
rect 38596 -6916 38624 -6908
rect 38632 -6916 38652 -6908
rect 38688 -6908 38772 -6888
rect 38688 -6916 38708 -6908
rect 38716 -6916 38744 -6908
rect 38752 -6916 38772 -6908
rect 38808 -6908 38892 -6888
rect 38808 -6916 38828 -6908
rect 38836 -6916 38864 -6908
rect 38872 -6916 38892 -6908
rect 38928 -6908 39012 -6888
rect 38928 -6916 38948 -6908
rect 38956 -6916 38984 -6908
rect 38992 -6916 39012 -6908
rect 39048 -6908 39132 -6888
rect 39048 -6916 39068 -6908
rect 39076 -6916 39104 -6908
rect 39112 -6916 39132 -6908
rect 39168 -6908 39252 -6888
rect 39168 -6916 39188 -6908
rect 39196 -6916 39224 -6908
rect 39232 -6916 39252 -6908
rect 39288 -6908 39372 -6888
rect 39288 -6916 39308 -6908
rect 39316 -6916 39344 -6908
rect 39352 -6916 39372 -6908
rect 39408 -6908 39492 -6888
rect 39408 -6916 39428 -6908
rect 39436 -6916 39464 -6908
rect 39472 -6916 39492 -6908
rect 39528 -6908 39612 -6888
rect 39528 -6916 39548 -6908
rect 39556 -6916 39584 -6908
rect 39592 -6916 39612 -6908
rect 39648 -6908 39732 -6888
rect 39648 -6916 39668 -6908
rect 39676 -6916 39704 -6908
rect 39712 -6916 39732 -6908
rect 39768 -6908 39852 -6888
rect 39768 -6916 39788 -6908
rect 39796 -6916 39824 -6908
rect 39832 -6916 39852 -6908
rect 39888 -6908 39972 -6888
rect 39888 -6916 39908 -6908
rect 39916 -6916 39944 -6908
rect 39952 -6916 39972 -6908
rect 40008 -6908 40092 -6888
rect 40008 -6916 40028 -6908
rect 40036 -6916 40064 -6908
rect 40072 -6916 40092 -6908
rect 40128 -6908 40212 -6888
rect 40128 -6916 40148 -6908
rect 40156 -6916 40184 -6908
rect 40192 -6916 40212 -6908
rect 40248 -6908 40332 -6888
rect 40248 -6916 40268 -6908
rect 40276 -6916 40304 -6908
rect 40312 -6916 40332 -6908
rect 40368 -6908 40452 -6888
rect 40368 -6916 40388 -6908
rect 40396 -6916 40424 -6908
rect 40432 -6916 40452 -6908
rect 40488 -6908 40572 -6888
rect 40488 -6916 40508 -6908
rect 40516 -6916 40544 -6908
rect 40552 -6916 40572 -6908
rect 40608 -6908 40692 -6888
rect 40608 -6916 40628 -6908
rect 40636 -6916 40664 -6908
rect 40672 -6916 40692 -6908
rect 40728 -6908 40812 -6888
rect 40728 -6916 40748 -6908
rect 40756 -6916 40784 -6908
rect 40792 -6916 40812 -6908
rect 40848 -6908 40932 -6888
rect 40848 -6916 40868 -6908
rect 40876 -6916 40904 -6908
rect 40912 -6916 40932 -6908
rect 40968 -6908 41052 -6888
rect 40968 -6916 40988 -6908
rect 40996 -6916 41024 -6908
rect 41032 -6916 41052 -6908
rect 41088 -6908 41172 -6888
rect 41088 -6916 41108 -6908
rect 41116 -6916 41144 -6908
rect 41152 -6916 41172 -6908
rect 41208 -6908 41292 -6888
rect 41208 -6916 41228 -6908
rect 41236 -6916 41264 -6908
rect 41272 -6916 41292 -6908
rect 41328 -6908 41412 -6888
rect 41328 -6916 41348 -6908
rect 41356 -6916 41384 -6908
rect 41392 -6916 41412 -6908
rect 41448 -6908 41532 -6888
rect 41448 -6916 41468 -6908
rect 41476 -6916 41504 -6908
rect 41512 -6916 41532 -6908
rect 41568 -6908 41652 -6888
rect 41568 -6916 41588 -6908
rect 41596 -6916 41624 -6908
rect 41632 -6916 41652 -6908
rect 41688 -6908 41772 -6888
rect 41688 -6916 41708 -6908
rect 41716 -6916 41744 -6908
rect 41752 -6916 41772 -6908
rect 41808 -6908 41892 -6888
rect 41808 -6916 41828 -6908
rect 41836 -6916 41864 -6908
rect 41872 -6916 41892 -6908
rect 41928 -6908 42012 -6888
rect 41928 -6916 41948 -6908
rect 41956 -6916 41984 -6908
rect 41992 -6916 42012 -6908
rect 42048 -6908 42132 -6888
rect 42048 -6916 42068 -6908
rect 42076 -6916 42104 -6908
rect 42112 -6916 42132 -6908
rect 42168 -6908 42252 -6888
rect 42168 -6916 42188 -6908
rect 42196 -6916 42224 -6908
rect 42232 -6916 42252 -6908
rect 42288 -6908 42372 -6888
rect 42288 -6916 42308 -6908
rect 42316 -6916 42344 -6908
rect 42352 -6916 42372 -6908
rect 42408 -6908 42492 -6888
rect 42408 -6916 42428 -6908
rect 42436 -6916 42464 -6908
rect 42472 -6916 42492 -6908
rect 42528 -6908 42612 -6888
rect 42528 -6916 42548 -6908
rect 42556 -6916 42584 -6908
rect 42592 -6916 42612 -6908
rect 42648 -6908 42732 -6888
rect 42648 -6916 42668 -6908
rect 42676 -6916 42704 -6908
rect 42712 -6916 42732 -6908
rect 42768 -6908 42852 -6888
rect 42768 -6916 42788 -6908
rect 42796 -6916 42824 -6908
rect 42832 -6916 42852 -6908
rect 42888 -6908 42972 -6888
rect 42888 -6916 42908 -6908
rect 42916 -6916 42944 -6908
rect 42952 -6916 42972 -6908
rect 43008 -6908 43092 -6888
rect 43008 -6916 43028 -6908
rect 43036 -6916 43064 -6908
rect 43072 -6916 43092 -6908
rect 43128 -6908 43212 -6888
rect 43128 -6916 43148 -6908
rect 43156 -6916 43184 -6908
rect 43192 -6916 43212 -6908
rect 43248 -6908 43332 -6888
rect 43248 -6916 43268 -6908
rect 43276 -6916 43304 -6908
rect 43312 -6916 43332 -6908
rect 43368 -6908 43452 -6888
rect 43368 -6916 43388 -6908
rect 43396 -6916 43424 -6908
rect 43432 -6916 43452 -6908
rect 43488 -6908 43572 -6888
rect 43488 -6916 43508 -6908
rect 43516 -6916 43544 -6908
rect 43552 -6916 43572 -6908
rect 43608 -6908 43692 -6888
rect 43608 -6916 43628 -6908
rect 43636 -6916 43664 -6908
rect 43672 -6916 43692 -6908
rect 43728 -6908 43812 -6888
rect 43728 -6916 43748 -6908
rect 43756 -6916 43784 -6908
rect 43792 -6916 43812 -6908
rect 43848 -6908 43932 -6888
rect 43848 -6916 43868 -6908
rect 43876 -6916 43904 -6908
rect 43912 -6916 43932 -6908
rect 43968 -6908 44052 -6888
rect 43968 -6916 43988 -6908
rect 43996 -6916 44024 -6908
rect 44032 -6916 44052 -6908
rect 44088 -6908 44172 -6888
rect 44088 -6916 44108 -6908
rect 44116 -6916 44144 -6908
rect 44152 -6916 44172 -6908
rect 44208 -6908 44292 -6888
rect 44208 -6916 44228 -6908
rect 44236 -6916 44264 -6908
rect 44272 -6916 44292 -6908
rect 44328 -6908 44412 -6888
rect 44328 -6916 44348 -6908
rect 44356 -6916 44384 -6908
rect 44392 -6916 44412 -6908
rect 44448 -6908 44532 -6888
rect 44448 -6916 44468 -6908
rect 44476 -6916 44504 -6908
rect 44512 -6916 44532 -6908
rect 44568 -6908 44652 -6888
rect 44568 -6916 44588 -6908
rect 44596 -6916 44624 -6908
rect 44632 -6916 44652 -6908
rect 44688 -6908 44772 -6888
rect 44688 -6916 44708 -6908
rect 44716 -6916 44744 -6908
rect 44752 -6916 44772 -6908
rect 44808 -6908 44892 -6888
rect 44808 -6916 44828 -6908
rect 44836 -6916 44864 -6908
rect 44872 -6916 44892 -6908
rect 44928 -6908 45012 -6888
rect 44928 -6916 44948 -6908
rect 44956 -6916 44984 -6908
rect 44992 -6916 45012 -6908
rect 45048 -6908 45132 -6888
rect 45048 -6916 45068 -6908
rect 45076 -6916 45104 -6908
rect 45112 -6916 45132 -6908
rect 45168 -6908 45252 -6888
rect 45168 -6916 45188 -6908
rect 45196 -6916 45224 -6908
rect 45232 -6916 45252 -6908
rect 45288 -6908 45372 -6888
rect 45288 -6916 45308 -6908
rect 45316 -6916 45344 -6908
rect 45352 -6916 45372 -6908
rect 45408 -6908 45492 -6888
rect 45408 -6916 45428 -6908
rect 45436 -6916 45464 -6908
rect 45472 -6916 45492 -6908
rect 45528 -6908 45612 -6888
rect 45528 -6916 45548 -6908
rect 45556 -6916 45584 -6908
rect 45592 -6916 45612 -6908
rect 25876 -6944 25932 -6916
rect 25996 -6944 26052 -6916
rect 26116 -6944 26172 -6916
rect 26236 -6944 26292 -6916
rect 26356 -6944 26412 -6916
rect 26476 -6944 26532 -6916
rect 26596 -6944 26652 -6916
rect 26716 -6944 26772 -6916
rect 26836 -6944 26892 -6916
rect 26956 -6944 27012 -6916
rect 27076 -6944 27132 -6916
rect 27196 -6944 27252 -6916
rect 27316 -6944 27372 -6916
rect 27436 -6944 27492 -6916
rect 27556 -6944 27612 -6916
rect 27676 -6944 27732 -6916
rect 27796 -6944 27852 -6916
rect 27916 -6944 27972 -6916
rect 28036 -6944 28092 -6916
rect 28156 -6944 28212 -6916
rect 28276 -6944 28332 -6916
rect 28396 -6944 28452 -6916
rect 28516 -6944 28572 -6916
rect 28636 -6944 28692 -6916
rect 28756 -6944 28812 -6916
rect 28876 -6944 28932 -6916
rect 28996 -6944 29052 -6916
rect 29116 -6944 29172 -6916
rect 29236 -6944 29292 -6916
rect 29356 -6944 29412 -6916
rect 29476 -6944 29532 -6916
rect 29596 -6944 29652 -6916
rect 29716 -6944 29772 -6916
rect 29836 -6944 29892 -6916
rect 29956 -6944 30012 -6916
rect 30076 -6944 30132 -6916
rect 30196 -6944 30252 -6916
rect 30316 -6944 30372 -6916
rect 30436 -6944 30492 -6916
rect 30556 -6944 30612 -6916
rect 30676 -6944 30732 -6916
rect 30796 -6944 30852 -6916
rect 30916 -6944 30972 -6916
rect 31036 -6944 31092 -6916
rect 31156 -6944 31212 -6916
rect 31276 -6944 31332 -6916
rect 31396 -6944 31452 -6916
rect 31516 -6944 31572 -6916
rect 31636 -6944 31692 -6916
rect 31756 -6944 31812 -6916
rect 31876 -6944 31932 -6916
rect 31996 -6944 32052 -6916
rect 32116 -6944 32172 -6916
rect 32236 -6944 32292 -6916
rect 32356 -6944 32412 -6916
rect 32476 -6944 32532 -6916
rect 32596 -6944 32652 -6916
rect 32716 -6944 32772 -6916
rect 32836 -6944 32892 -6916
rect 32956 -6944 33012 -6916
rect 33076 -6944 33132 -6916
rect 33196 -6944 33252 -6916
rect 33316 -6944 33372 -6916
rect 33436 -6944 33492 -6916
rect 33556 -6944 33612 -6916
rect 33676 -6944 33732 -6916
rect 33796 -6944 33852 -6916
rect 33916 -6944 33972 -6916
rect 34036 -6944 34092 -6916
rect 34156 -6944 34212 -6916
rect 34276 -6944 34332 -6916
rect 34396 -6944 34452 -6916
rect 34516 -6944 34572 -6916
rect 34636 -6944 34692 -6916
rect 34756 -6944 34812 -6916
rect 34876 -6944 34932 -6916
rect 34996 -6944 35052 -6916
rect 35116 -6944 35172 -6916
rect 35236 -6944 35292 -6916
rect 35356 -6944 35412 -6916
rect 35476 -6944 35532 -6916
rect 35596 -6944 35652 -6916
rect 35716 -6944 35772 -6916
rect 35836 -6944 35892 -6916
rect 35956 -6944 36012 -6916
rect 36076 -6944 36132 -6916
rect 36196 -6944 36252 -6916
rect 36316 -6944 36372 -6916
rect 36436 -6944 36492 -6916
rect 36556 -6944 36612 -6916
rect 36676 -6944 36732 -6916
rect 36796 -6944 36852 -6916
rect 36916 -6944 36972 -6916
rect 37036 -6944 37092 -6916
rect 37156 -6944 37212 -6916
rect 37276 -6944 37332 -6916
rect 37396 -6944 37452 -6916
rect 37516 -6944 37572 -6916
rect 37636 -6944 37692 -6916
rect 37756 -6944 37812 -6916
rect 37876 -6944 37932 -6916
rect 37996 -6944 38052 -6916
rect 38116 -6944 38172 -6916
rect 38236 -6944 38292 -6916
rect 38356 -6944 38412 -6916
rect 38476 -6944 38532 -6916
rect 38596 -6944 38652 -6916
rect 38716 -6944 38772 -6916
rect 38836 -6944 38892 -6916
rect 38956 -6944 39012 -6916
rect 39076 -6944 39132 -6916
rect 39196 -6944 39252 -6916
rect 39316 -6944 39372 -6916
rect 39436 -6944 39492 -6916
rect 39556 -6944 39612 -6916
rect 39676 -6944 39732 -6916
rect 39796 -6944 39852 -6916
rect 39916 -6944 39972 -6916
rect 40036 -6944 40092 -6916
rect 40156 -6944 40212 -6916
rect 40276 -6944 40332 -6916
rect 40396 -6944 40452 -6916
rect 40516 -6944 40572 -6916
rect 40636 -6944 40692 -6916
rect 40756 -6944 40812 -6916
rect 40876 -6944 40932 -6916
rect 40996 -6944 41052 -6916
rect 41116 -6944 41172 -6916
rect 41236 -6944 41292 -6916
rect 41356 -6944 41412 -6916
rect 41476 -6944 41532 -6916
rect 41596 -6944 41652 -6916
rect 41716 -6944 41772 -6916
rect 41836 -6944 41892 -6916
rect 41956 -6944 42012 -6916
rect 42076 -6944 42132 -6916
rect 42196 -6944 42252 -6916
rect 42316 -6944 42372 -6916
rect 42436 -6944 42492 -6916
rect 42556 -6944 42612 -6916
rect 42676 -6944 42732 -6916
rect 42796 -6944 42852 -6916
rect 42916 -6944 42972 -6916
rect 43036 -6944 43092 -6916
rect 43156 -6944 43212 -6916
rect 43276 -6944 43332 -6916
rect 43396 -6944 43452 -6916
rect 43516 -6944 43572 -6916
rect 43636 -6944 43692 -6916
rect 43756 -6944 43812 -6916
rect 43876 -6944 43932 -6916
rect 43996 -6944 44052 -6916
rect 44116 -6944 44172 -6916
rect 44236 -6944 44292 -6916
rect 44356 -6944 44412 -6916
rect 44476 -6944 44532 -6916
rect 44596 -6944 44652 -6916
rect 44716 -6944 44772 -6916
rect 44836 -6944 44892 -6916
rect 44956 -6944 45012 -6916
rect 45076 -6944 45132 -6916
rect 45196 -6944 45252 -6916
rect 45316 -6944 45372 -6916
rect 45436 -6944 45492 -6916
rect 45556 -6944 45612 -6916
rect 25848 -12008 25932 -11988
rect 25848 -12016 25868 -12008
rect 25876 -12016 25904 -12008
rect 25912 -12016 25932 -12008
rect 26088 -12008 26172 -11988
rect 26088 -12016 26108 -12008
rect 26116 -12016 26144 -12008
rect 26152 -12016 26172 -12008
rect 26208 -12008 26292 -11988
rect 26208 -12016 26228 -12008
rect 26236 -12016 26264 -12008
rect 26272 -12016 26292 -12008
rect 26448 -12008 26532 -11988
rect 26448 -12016 26468 -12008
rect 26476 -12016 26504 -12008
rect 26512 -12016 26532 -12008
rect 26568 -12008 26652 -11988
rect 26568 -12016 26588 -12008
rect 26596 -12016 26624 -12008
rect 26632 -12016 26652 -12008
rect 26808 -12008 26892 -11988
rect 26808 -12016 26828 -12008
rect 26836 -12016 26864 -12008
rect 26872 -12016 26892 -12008
rect 26928 -12008 27012 -11988
rect 26928 -12016 26948 -12008
rect 26956 -12016 26984 -12008
rect 26992 -12016 27012 -12008
rect 27168 -12008 27252 -11988
rect 27168 -12016 27188 -12008
rect 27196 -12016 27224 -12008
rect 27232 -12016 27252 -12008
rect 27288 -12008 27372 -11988
rect 27288 -12016 27308 -12008
rect 27316 -12016 27344 -12008
rect 27352 -12016 27372 -12008
rect 27528 -12008 27612 -11988
rect 27528 -12016 27548 -12008
rect 27556 -12016 27584 -12008
rect 27592 -12016 27612 -12008
rect 27648 -12008 27732 -11988
rect 27648 -12016 27668 -12008
rect 27676 -12016 27704 -12008
rect 27712 -12016 27732 -12008
rect 27888 -12008 27972 -11988
rect 27888 -12016 27908 -12008
rect 27916 -12016 27944 -12008
rect 27952 -12016 27972 -12008
rect 28008 -12008 28092 -11988
rect 28008 -12016 28028 -12008
rect 28036 -12016 28064 -12008
rect 28072 -12016 28092 -12008
rect 28248 -12008 28332 -11988
rect 28248 -12016 28268 -12008
rect 28276 -12016 28304 -12008
rect 28312 -12016 28332 -12008
rect 28368 -12008 28452 -11988
rect 28368 -12016 28388 -12008
rect 28396 -12016 28424 -12008
rect 28432 -12016 28452 -12008
rect 28608 -12008 28692 -11988
rect 28608 -12016 28628 -12008
rect 28636 -12016 28664 -12008
rect 28672 -12016 28692 -12008
rect 28728 -12008 28812 -11988
rect 28728 -12016 28748 -12008
rect 28756 -12016 28784 -12008
rect 28792 -12016 28812 -12008
rect 28968 -12008 29052 -11988
rect 28968 -12016 28988 -12008
rect 28996 -12016 29024 -12008
rect 29032 -12016 29052 -12008
rect 29088 -12008 29172 -11988
rect 29088 -12016 29108 -12008
rect 29116 -12016 29144 -12008
rect 29152 -12016 29172 -12008
rect 29328 -12008 29412 -11988
rect 29328 -12016 29348 -12008
rect 29356 -12016 29384 -12008
rect 29392 -12016 29412 -12008
rect 29448 -12008 29532 -11988
rect 29448 -12016 29468 -12008
rect 29476 -12016 29504 -12008
rect 29512 -12016 29532 -12008
rect 29688 -12008 29772 -11988
rect 29688 -12016 29708 -12008
rect 29716 -12016 29744 -12008
rect 29752 -12016 29772 -12008
rect 29808 -12008 29892 -11988
rect 29808 -12016 29828 -12008
rect 29836 -12016 29864 -12008
rect 29872 -12016 29892 -12008
rect 30048 -12008 30132 -11988
rect 30048 -12016 30068 -12008
rect 30076 -12016 30104 -12008
rect 30112 -12016 30132 -12008
rect 30168 -12008 30252 -11988
rect 30168 -12016 30188 -12008
rect 30196 -12016 30224 -12008
rect 30232 -12016 30252 -12008
rect 30408 -12008 30492 -11988
rect 30408 -12016 30428 -12008
rect 30436 -12016 30464 -12008
rect 30472 -12016 30492 -12008
rect 30528 -12008 30612 -11988
rect 30528 -12016 30548 -12008
rect 30556 -12016 30584 -12008
rect 30592 -12016 30612 -12008
rect 30768 -12008 30852 -11988
rect 30768 -12016 30788 -12008
rect 30796 -12016 30824 -12008
rect 30832 -12016 30852 -12008
rect 30888 -12008 30972 -11988
rect 30888 -12016 30908 -12008
rect 30916 -12016 30944 -12008
rect 30952 -12016 30972 -12008
rect 31128 -12008 31212 -11988
rect 31128 -12016 31148 -12008
rect 31156 -12016 31184 -12008
rect 31192 -12016 31212 -12008
rect 31248 -12008 31332 -11988
rect 31248 -12016 31268 -12008
rect 31276 -12016 31304 -12008
rect 31312 -12016 31332 -12008
rect 31488 -12008 31572 -11988
rect 31488 -12016 31508 -12008
rect 31516 -12016 31544 -12008
rect 31552 -12016 31572 -12008
rect 31608 -12008 31692 -11988
rect 31608 -12016 31628 -12008
rect 31636 -12016 31664 -12008
rect 31672 -12016 31692 -12008
rect 31848 -12008 31932 -11988
rect 31848 -12016 31868 -12008
rect 31876 -12016 31904 -12008
rect 31912 -12016 31932 -12008
rect 31968 -12008 32052 -11988
rect 31968 -12016 31988 -12008
rect 31996 -12016 32024 -12008
rect 32032 -12016 32052 -12008
rect 32208 -12008 32292 -11988
rect 32208 -12016 32228 -12008
rect 32236 -12016 32264 -12008
rect 32272 -12016 32292 -12008
rect 32328 -12008 32412 -11988
rect 32328 -12016 32348 -12008
rect 32356 -12016 32384 -12008
rect 32392 -12016 32412 -12008
rect 32568 -12008 32652 -11988
rect 32568 -12016 32588 -12008
rect 32596 -12016 32624 -12008
rect 32632 -12016 32652 -12008
rect 32688 -12008 32772 -11988
rect 32688 -12016 32708 -12008
rect 32716 -12016 32744 -12008
rect 32752 -12016 32772 -12008
rect 32928 -12008 33012 -11988
rect 32928 -12016 32948 -12008
rect 32956 -12016 32984 -12008
rect 32992 -12016 33012 -12008
rect 33048 -12008 33132 -11988
rect 33048 -12016 33068 -12008
rect 33076 -12016 33104 -12008
rect 33112 -12016 33132 -12008
rect 33288 -12008 33372 -11988
rect 33288 -12016 33308 -12008
rect 33316 -12016 33344 -12008
rect 33352 -12016 33372 -12008
rect 33408 -12008 33492 -11988
rect 33408 -12016 33428 -12008
rect 33436 -12016 33464 -12008
rect 33472 -12016 33492 -12008
rect 33648 -12008 33732 -11988
rect 33648 -12016 33668 -12008
rect 33676 -12016 33704 -12008
rect 33712 -12016 33732 -12008
rect 33768 -12008 33852 -11988
rect 33768 -12016 33788 -12008
rect 33796 -12016 33824 -12008
rect 33832 -12016 33852 -12008
rect 34008 -12008 34092 -11988
rect 34008 -12016 34028 -12008
rect 34036 -12016 34064 -12008
rect 34072 -12016 34092 -12008
rect 34128 -12008 34212 -11988
rect 34128 -12016 34148 -12008
rect 34156 -12016 34184 -12008
rect 34192 -12016 34212 -12008
rect 34368 -12008 34452 -11988
rect 34368 -12016 34388 -12008
rect 34396 -12016 34424 -12008
rect 34432 -12016 34452 -12008
rect 34488 -12008 34572 -11988
rect 34488 -12016 34508 -12008
rect 34516 -12016 34544 -12008
rect 34552 -12016 34572 -12008
rect 34728 -12008 34812 -11988
rect 34728 -12016 34748 -12008
rect 34756 -12016 34784 -12008
rect 34792 -12016 34812 -12008
rect 34848 -12008 34932 -11988
rect 34848 -12016 34868 -12008
rect 34876 -12016 34904 -12008
rect 34912 -12016 34932 -12008
rect 35088 -12008 35172 -11988
rect 35088 -12016 35108 -12008
rect 35116 -12016 35144 -12008
rect 35152 -12016 35172 -12008
rect 35208 -12008 35292 -11988
rect 35208 -12016 35228 -12008
rect 35236 -12016 35264 -12008
rect 35272 -12016 35292 -12008
rect 35448 -12008 35532 -11988
rect 35448 -12016 35468 -12008
rect 35476 -12016 35504 -12008
rect 35512 -12016 35532 -12008
rect 35568 -12008 35652 -11988
rect 35568 -12016 35588 -12008
rect 35596 -12016 35624 -12008
rect 35632 -12016 35652 -12008
rect 35808 -12008 35892 -11988
rect 35808 -12016 35828 -12008
rect 35836 -12016 35864 -12008
rect 35872 -12016 35892 -12008
rect 35928 -12008 36012 -11988
rect 35928 -12016 35948 -12008
rect 35956 -12016 35984 -12008
rect 35992 -12016 36012 -12008
rect 36168 -12008 36252 -11988
rect 36168 -12016 36188 -12008
rect 36196 -12016 36224 -12008
rect 36232 -12016 36252 -12008
rect 36288 -12008 36372 -11988
rect 36288 -12016 36308 -12008
rect 36316 -12016 36344 -12008
rect 36352 -12016 36372 -12008
rect 36528 -12008 36612 -11988
rect 36528 -12016 36548 -12008
rect 36556 -12016 36584 -12008
rect 36592 -12016 36612 -12008
rect 36648 -12008 36732 -11988
rect 36648 -12016 36668 -12008
rect 36676 -12016 36704 -12008
rect 36712 -12016 36732 -12008
rect 36888 -12008 36972 -11988
rect 36888 -12016 36908 -12008
rect 36916 -12016 36944 -12008
rect 36952 -12016 36972 -12008
rect 37008 -12008 37092 -11988
rect 37008 -12016 37028 -12008
rect 37036 -12016 37064 -12008
rect 37072 -12016 37092 -12008
rect 37248 -12008 37332 -11988
rect 37248 -12016 37268 -12008
rect 37276 -12016 37304 -12008
rect 37312 -12016 37332 -12008
rect 37368 -12008 37452 -11988
rect 37368 -12016 37388 -12008
rect 37396 -12016 37424 -12008
rect 37432 -12016 37452 -12008
rect 37608 -12008 37692 -11988
rect 37608 -12016 37628 -12008
rect 37636 -12016 37664 -12008
rect 37672 -12016 37692 -12008
rect 37728 -12008 37812 -11988
rect 37728 -12016 37748 -12008
rect 37756 -12016 37784 -12008
rect 37792 -12016 37812 -12008
rect 37968 -12008 38052 -11988
rect 37968 -12016 37988 -12008
rect 37996 -12016 38024 -12008
rect 38032 -12016 38052 -12008
rect 38088 -12008 38172 -11988
rect 38088 -12016 38108 -12008
rect 38116 -12016 38144 -12008
rect 38152 -12016 38172 -12008
rect 38328 -12008 38412 -11988
rect 38328 -12016 38348 -12008
rect 38356 -12016 38384 -12008
rect 38392 -12016 38412 -12008
rect 38448 -12008 38532 -11988
rect 38448 -12016 38468 -12008
rect 38476 -12016 38504 -12008
rect 38512 -12016 38532 -12008
rect 38688 -12008 38772 -11988
rect 38688 -12016 38708 -12008
rect 38716 -12016 38744 -12008
rect 38752 -12016 38772 -12008
rect 38808 -12008 38892 -11988
rect 38808 -12016 38828 -12008
rect 38836 -12016 38864 -12008
rect 38872 -12016 38892 -12008
rect 39048 -12008 39132 -11988
rect 39048 -12016 39068 -12008
rect 39076 -12016 39104 -12008
rect 39112 -12016 39132 -12008
rect 39168 -12008 39252 -11988
rect 39168 -12016 39188 -12008
rect 39196 -12016 39224 -12008
rect 39232 -12016 39252 -12008
rect 39408 -12008 39492 -11988
rect 39408 -12016 39428 -12008
rect 39436 -12016 39464 -12008
rect 39472 -12016 39492 -12008
rect 39528 -12008 39612 -11988
rect 39528 -12016 39548 -12008
rect 39556 -12016 39584 -12008
rect 39592 -12016 39612 -12008
rect 39768 -12008 39852 -11988
rect 39768 -12016 39788 -12008
rect 39796 -12016 39824 -12008
rect 39832 -12016 39852 -12008
rect 39888 -12008 39972 -11988
rect 39888 -12016 39908 -12008
rect 39916 -12016 39944 -12008
rect 39952 -12016 39972 -12008
rect 40128 -12008 40212 -11988
rect 40128 -12016 40148 -12008
rect 40156 -12016 40184 -12008
rect 40192 -12016 40212 -12008
rect 40248 -12008 40332 -11988
rect 40248 -12016 40268 -12008
rect 40276 -12016 40304 -12008
rect 40312 -12016 40332 -12008
rect 40488 -12008 40572 -11988
rect 40488 -12016 40508 -12008
rect 40516 -12016 40544 -12008
rect 40552 -12016 40572 -12008
rect 40608 -12008 40692 -11988
rect 40608 -12016 40628 -12008
rect 40636 -12016 40664 -12008
rect 40672 -12016 40692 -12008
rect 40848 -12008 40932 -11988
rect 40848 -12016 40868 -12008
rect 40876 -12016 40904 -12008
rect 40912 -12016 40932 -12008
rect 40968 -12008 41052 -11988
rect 40968 -12016 40988 -12008
rect 40996 -12016 41024 -12008
rect 41032 -12016 41052 -12008
rect 41208 -12008 41292 -11988
rect 41208 -12016 41228 -12008
rect 41236 -12016 41264 -12008
rect 41272 -12016 41292 -12008
rect 41328 -12008 41412 -11988
rect 41328 -12016 41348 -12008
rect 41356 -12016 41384 -12008
rect 41392 -12016 41412 -12008
rect 41568 -12008 41652 -11988
rect 41568 -12016 41588 -12008
rect 41596 -12016 41624 -12008
rect 41632 -12016 41652 -12008
rect 41688 -12008 41772 -11988
rect 41688 -12016 41708 -12008
rect 41716 -12016 41744 -12008
rect 41752 -12016 41772 -12008
rect 41928 -12008 42012 -11988
rect 41928 -12016 41948 -12008
rect 41956 -12016 41984 -12008
rect 41992 -12016 42012 -12008
rect 42048 -12008 42132 -11988
rect 42048 -12016 42068 -12008
rect 42076 -12016 42104 -12008
rect 42112 -12016 42132 -12008
rect 42288 -12008 42372 -11988
rect 42288 -12016 42308 -12008
rect 42316 -12016 42344 -12008
rect 42352 -12016 42372 -12008
rect 42408 -12008 42492 -11988
rect 42408 -12016 42428 -12008
rect 42436 -12016 42464 -12008
rect 42472 -12016 42492 -12008
rect 42648 -12008 42732 -11988
rect 42648 -12016 42668 -12008
rect 42676 -12016 42704 -12008
rect 42712 -12016 42732 -12008
rect 42768 -12008 42852 -11988
rect 42768 -12016 42788 -12008
rect 42796 -12016 42824 -12008
rect 42832 -12016 42852 -12008
rect 43008 -12008 43092 -11988
rect 43008 -12016 43028 -12008
rect 43036 -12016 43064 -12008
rect 43072 -12016 43092 -12008
rect 43128 -12008 43212 -11988
rect 43128 -12016 43148 -12008
rect 43156 -12016 43184 -12008
rect 43192 -12016 43212 -12008
rect 43248 -12008 43332 -11988
rect 43248 -12016 43268 -12008
rect 43276 -12016 43304 -12008
rect 43312 -12016 43332 -12008
rect 43488 -12008 43572 -11988
rect 43488 -12016 43508 -12008
rect 43516 -12016 43544 -12008
rect 43552 -12016 43572 -12008
rect 43608 -12008 43692 -11988
rect 43608 -12016 43628 -12008
rect 43636 -12016 43664 -12008
rect 43672 -12016 43692 -12008
rect 43848 -12008 43932 -11988
rect 43848 -12016 43868 -12008
rect 43876 -12016 43904 -12008
rect 43912 -12016 43932 -12008
rect 43968 -12008 44052 -11988
rect 43968 -12016 43988 -12008
rect 43996 -12016 44024 -12008
rect 44032 -12016 44052 -12008
rect 44208 -12008 44292 -11988
rect 44208 -12016 44228 -12008
rect 44236 -12016 44264 -12008
rect 44272 -12016 44292 -12008
rect 44328 -12008 44412 -11988
rect 44328 -12016 44348 -12008
rect 44356 -12016 44384 -12008
rect 44392 -12016 44412 -12008
rect 44448 -12008 44532 -11988
rect 44448 -12016 44468 -12008
rect 44476 -12016 44504 -12008
rect 44512 -12016 44532 -12008
rect 44688 -12008 44772 -11988
rect 44688 -12016 44708 -12008
rect 44716 -12016 44744 -12008
rect 44752 -12016 44772 -12008
rect 44808 -12008 44892 -11988
rect 44808 -12016 44828 -12008
rect 44836 -12016 44864 -12008
rect 44872 -12016 44892 -12008
rect 45048 -12008 45132 -11988
rect 45048 -12016 45068 -12008
rect 45076 -12016 45104 -12008
rect 45112 -12016 45132 -12008
rect 45168 -12008 45252 -11988
rect 45168 -12016 45188 -12008
rect 45196 -12016 45224 -12008
rect 45232 -12016 45252 -12008
rect 45408 -12008 45492 -11988
rect 45408 -12016 45428 -12008
rect 45436 -12016 45464 -12008
rect 45472 -12016 45492 -12008
rect 45528 -12008 45612 -11988
rect 45528 -12016 45548 -12008
rect 45556 -12016 45584 -12008
rect 45592 -12016 45612 -12008
rect 25876 -12044 25932 -12016
rect 26116 -12044 26172 -12016
rect 26236 -12044 26292 -12016
rect 26476 -12044 26532 -12016
rect 26596 -12044 26652 -12016
rect 26836 -12044 26892 -12016
rect 26956 -12044 27012 -12016
rect 27196 -12044 27252 -12016
rect 27316 -12044 27372 -12016
rect 27556 -12044 27612 -12016
rect 27676 -12044 27732 -12016
rect 27916 -12044 27972 -12016
rect 28036 -12044 28092 -12016
rect 28276 -12044 28332 -12016
rect 28396 -12044 28452 -12016
rect 28636 -12044 28692 -12016
rect 28756 -12044 28812 -12016
rect 28996 -12044 29052 -12016
rect 29116 -12044 29172 -12016
rect 29356 -12044 29412 -12016
rect 29476 -12044 29532 -12016
rect 29716 -12044 29772 -12016
rect 29836 -12044 29892 -12016
rect 30076 -12044 30132 -12016
rect 30196 -12044 30252 -12016
rect 30436 -12044 30492 -12016
rect 30556 -12044 30612 -12016
rect 30796 -12044 30852 -12016
rect 30916 -12044 30972 -12016
rect 31156 -12044 31212 -12016
rect 31276 -12044 31332 -12016
rect 31516 -12044 31572 -12016
rect 31636 -12044 31692 -12016
rect 31876 -12044 31932 -12016
rect 31996 -12044 32052 -12016
rect 32236 -12044 32292 -12016
rect 32356 -12044 32412 -12016
rect 32596 -12044 32652 -12016
rect 32716 -12044 32772 -12016
rect 32956 -12044 33012 -12016
rect 33076 -12044 33132 -12016
rect 33316 -12044 33372 -12016
rect 33436 -12044 33492 -12016
rect 33676 -12044 33732 -12016
rect 33796 -12044 33852 -12016
rect 34036 -12044 34092 -12016
rect 34156 -12044 34212 -12016
rect 34396 -12044 34452 -12016
rect 34516 -12044 34572 -12016
rect 34756 -12044 34812 -12016
rect 34876 -12044 34932 -12016
rect 35116 -12044 35172 -12016
rect 35236 -12044 35292 -12016
rect 35476 -12044 35532 -12016
rect 35596 -12044 35652 -12016
rect 35836 -12044 35892 -12016
rect 35956 -12044 36012 -12016
rect 36196 -12044 36252 -12016
rect 36316 -12044 36372 -12016
rect 36556 -12044 36612 -12016
rect 36676 -12044 36732 -12016
rect 36916 -12044 36972 -12016
rect 37036 -12044 37092 -12016
rect 37276 -12044 37332 -12016
rect 37396 -12044 37452 -12016
rect 37636 -12044 37692 -12016
rect 37756 -12044 37812 -12016
rect 37996 -12044 38052 -12016
rect 38116 -12044 38172 -12016
rect 38356 -12044 38412 -12016
rect 38476 -12044 38532 -12016
rect 38716 -12044 38772 -12016
rect 38836 -12044 38892 -12016
rect 39076 -12044 39132 -12016
rect 39196 -12044 39252 -12016
rect 39436 -12044 39492 -12016
rect 39556 -12044 39612 -12016
rect 39796 -12044 39852 -12016
rect 39916 -12044 39972 -12016
rect 40156 -12044 40212 -12016
rect 40276 -12044 40332 -12016
rect 40516 -12044 40572 -12016
rect 40636 -12044 40692 -12016
rect 40876 -12044 40932 -12016
rect 40996 -12044 41052 -12016
rect 41236 -12044 41292 -12016
rect 41356 -12044 41412 -12016
rect 41596 -12044 41652 -12016
rect 41716 -12044 41772 -12016
rect 41956 -12044 42012 -12016
rect 42076 -12044 42132 -12016
rect 42316 -12044 42372 -12016
rect 42436 -12044 42492 -12016
rect 42676 -12044 42732 -12016
rect 42796 -12044 42852 -12016
rect 43036 -12044 43092 -12016
rect 43156 -12044 43212 -12016
rect 43276 -12044 43332 -12016
rect 43516 -12044 43572 -12016
rect 43636 -12044 43692 -12016
rect 43876 -12044 43932 -12016
rect 43996 -12044 44052 -12016
rect 44236 -12044 44292 -12016
rect 44356 -12044 44412 -12016
rect 44476 -12044 44532 -12016
rect 44716 -12044 44772 -12016
rect 44836 -12044 44892 -12016
rect 45076 -12044 45132 -12016
rect 45196 -12044 45252 -12016
rect 45436 -12044 45492 -12016
rect 45556 -12044 45612 -12016
rect 25848 -12188 25932 -12168
rect 25848 -12196 25868 -12188
rect 25876 -12196 25904 -12188
rect 25912 -12196 25932 -12188
rect 25968 -12188 26052 -12168
rect 25968 -12196 25988 -12188
rect 25996 -12196 26024 -12188
rect 26032 -12196 26052 -12188
rect 26088 -12188 26172 -12168
rect 26088 -12196 26108 -12188
rect 26116 -12196 26144 -12188
rect 26152 -12196 26172 -12188
rect 26208 -12188 26292 -12168
rect 26208 -12196 26228 -12188
rect 26236 -12196 26264 -12188
rect 26272 -12196 26292 -12188
rect 26328 -12188 26412 -12168
rect 26328 -12196 26348 -12188
rect 26356 -12196 26384 -12188
rect 26392 -12196 26412 -12188
rect 26448 -12188 26532 -12168
rect 26448 -12196 26468 -12188
rect 26476 -12196 26504 -12188
rect 26512 -12196 26532 -12188
rect 26568 -12188 26652 -12168
rect 26568 -12196 26588 -12188
rect 26596 -12196 26624 -12188
rect 26632 -12196 26652 -12188
rect 26688 -12188 26772 -12168
rect 26688 -12196 26708 -12188
rect 26716 -12196 26744 -12188
rect 26752 -12196 26772 -12188
rect 26808 -12188 26892 -12168
rect 26808 -12196 26828 -12188
rect 26836 -12196 26864 -12188
rect 26872 -12196 26892 -12188
rect 26928 -12188 27012 -12168
rect 26928 -12196 26948 -12188
rect 26956 -12196 26984 -12188
rect 26992 -12196 27012 -12188
rect 27048 -12188 27132 -12168
rect 27048 -12196 27068 -12188
rect 27076 -12196 27104 -12188
rect 27112 -12196 27132 -12188
rect 27168 -12188 27252 -12168
rect 27168 -12196 27188 -12188
rect 27196 -12196 27224 -12188
rect 27232 -12196 27252 -12188
rect 27288 -12188 27372 -12168
rect 27288 -12196 27308 -12188
rect 27316 -12196 27344 -12188
rect 27352 -12196 27372 -12188
rect 27408 -12188 27492 -12168
rect 27408 -12196 27428 -12188
rect 27436 -12196 27464 -12188
rect 27472 -12196 27492 -12188
rect 27528 -12188 27612 -12168
rect 27528 -12196 27548 -12188
rect 27556 -12196 27584 -12188
rect 27592 -12196 27612 -12188
rect 27648 -12188 27732 -12168
rect 27648 -12196 27668 -12188
rect 27676 -12196 27704 -12188
rect 27712 -12196 27732 -12188
rect 27768 -12188 27852 -12168
rect 27768 -12196 27788 -12188
rect 27796 -12196 27824 -12188
rect 27832 -12196 27852 -12188
rect 27888 -12188 27972 -12168
rect 27888 -12196 27908 -12188
rect 27916 -12196 27944 -12188
rect 27952 -12196 27972 -12188
rect 28008 -12188 28092 -12168
rect 28008 -12196 28028 -12188
rect 28036 -12196 28064 -12188
rect 28072 -12196 28092 -12188
rect 28128 -12188 28212 -12168
rect 28128 -12196 28148 -12188
rect 28156 -12196 28184 -12188
rect 28192 -12196 28212 -12188
rect 28248 -12188 28332 -12168
rect 28248 -12196 28268 -12188
rect 28276 -12196 28304 -12188
rect 28312 -12196 28332 -12188
rect 28368 -12188 28452 -12168
rect 28368 -12196 28388 -12188
rect 28396 -12196 28424 -12188
rect 28432 -12196 28452 -12188
rect 28488 -12188 28572 -12168
rect 28488 -12196 28508 -12188
rect 28516 -12196 28544 -12188
rect 28552 -12196 28572 -12188
rect 28608 -12188 28692 -12168
rect 28608 -12196 28628 -12188
rect 28636 -12196 28664 -12188
rect 28672 -12196 28692 -12188
rect 28728 -12188 28812 -12168
rect 28728 -12196 28748 -12188
rect 28756 -12196 28784 -12188
rect 28792 -12196 28812 -12188
rect 28848 -12188 28932 -12168
rect 28848 -12196 28868 -12188
rect 28876 -12196 28904 -12188
rect 28912 -12196 28932 -12188
rect 28968 -12188 29052 -12168
rect 28968 -12196 28988 -12188
rect 28996 -12196 29024 -12188
rect 29032 -12196 29052 -12188
rect 29088 -12188 29172 -12168
rect 29088 -12196 29108 -12188
rect 29116 -12196 29144 -12188
rect 29152 -12196 29172 -12188
rect 29208 -12188 29292 -12168
rect 29208 -12196 29228 -12188
rect 29236 -12196 29264 -12188
rect 29272 -12196 29292 -12188
rect 29328 -12188 29412 -12168
rect 29328 -12196 29348 -12188
rect 29356 -12196 29384 -12188
rect 29392 -12196 29412 -12188
rect 29448 -12188 29532 -12168
rect 29448 -12196 29468 -12188
rect 29476 -12196 29504 -12188
rect 29512 -12196 29532 -12188
rect 29568 -12188 29652 -12168
rect 29568 -12196 29588 -12188
rect 29596 -12196 29624 -12188
rect 29632 -12196 29652 -12188
rect 29688 -12188 29772 -12168
rect 29688 -12196 29708 -12188
rect 29716 -12196 29744 -12188
rect 29752 -12196 29772 -12188
rect 29808 -12188 29892 -12168
rect 29808 -12196 29828 -12188
rect 29836 -12196 29864 -12188
rect 29872 -12196 29892 -12188
rect 29928 -12188 30012 -12168
rect 29928 -12196 29948 -12188
rect 29956 -12196 29984 -12188
rect 29992 -12196 30012 -12188
rect 30048 -12188 30132 -12168
rect 30048 -12196 30068 -12188
rect 30076 -12196 30104 -12188
rect 30112 -12196 30132 -12188
rect 30168 -12188 30252 -12168
rect 30168 -12196 30188 -12188
rect 30196 -12196 30224 -12188
rect 30232 -12196 30252 -12188
rect 30288 -12188 30372 -12168
rect 30288 -12196 30308 -12188
rect 30316 -12196 30344 -12188
rect 30352 -12196 30372 -12188
rect 30408 -12188 30492 -12168
rect 30408 -12196 30428 -12188
rect 30436 -12196 30464 -12188
rect 30472 -12196 30492 -12188
rect 30528 -12188 30612 -12168
rect 30528 -12196 30548 -12188
rect 30556 -12196 30584 -12188
rect 30592 -12196 30612 -12188
rect 30648 -12188 30732 -12168
rect 30648 -12196 30668 -12188
rect 30676 -12196 30704 -12188
rect 30712 -12196 30732 -12188
rect 30768 -12188 30852 -12168
rect 30768 -12196 30788 -12188
rect 30796 -12196 30824 -12188
rect 30832 -12196 30852 -12188
rect 30888 -12188 30972 -12168
rect 30888 -12196 30908 -12188
rect 30916 -12196 30944 -12188
rect 30952 -12196 30972 -12188
rect 31008 -12188 31092 -12168
rect 31008 -12196 31028 -12188
rect 31036 -12196 31064 -12188
rect 31072 -12196 31092 -12188
rect 31128 -12188 31212 -12168
rect 31128 -12196 31148 -12188
rect 31156 -12196 31184 -12188
rect 31192 -12196 31212 -12188
rect 31248 -12188 31332 -12168
rect 31248 -12196 31268 -12188
rect 31276 -12196 31304 -12188
rect 31312 -12196 31332 -12188
rect 31368 -12188 31452 -12168
rect 31368 -12196 31388 -12188
rect 31396 -12196 31424 -12188
rect 31432 -12196 31452 -12188
rect 31488 -12188 31572 -12168
rect 31488 -12196 31508 -12188
rect 31516 -12196 31544 -12188
rect 31552 -12196 31572 -12188
rect 31608 -12188 31692 -12168
rect 31608 -12196 31628 -12188
rect 31636 -12196 31664 -12188
rect 31672 -12196 31692 -12188
rect 31728 -12188 31812 -12168
rect 31728 -12196 31748 -12188
rect 31756 -12196 31784 -12188
rect 31792 -12196 31812 -12188
rect 31848 -12188 31932 -12168
rect 31848 -12196 31868 -12188
rect 31876 -12196 31904 -12188
rect 31912 -12196 31932 -12188
rect 31968 -12188 32052 -12168
rect 31968 -12196 31988 -12188
rect 31996 -12196 32024 -12188
rect 32032 -12196 32052 -12188
rect 32088 -12188 32172 -12168
rect 32088 -12196 32108 -12188
rect 32116 -12196 32144 -12188
rect 32152 -12196 32172 -12188
rect 32208 -12188 32292 -12168
rect 32208 -12196 32228 -12188
rect 32236 -12196 32264 -12188
rect 32272 -12196 32292 -12188
rect 32328 -12188 32412 -12168
rect 32328 -12196 32348 -12188
rect 32356 -12196 32384 -12188
rect 32392 -12196 32412 -12188
rect 32448 -12188 32532 -12168
rect 32448 -12196 32468 -12188
rect 32476 -12196 32504 -12188
rect 32512 -12196 32532 -12188
rect 32568 -12188 32652 -12168
rect 32568 -12196 32588 -12188
rect 32596 -12196 32624 -12188
rect 32632 -12196 32652 -12188
rect 32688 -12188 32772 -12168
rect 32688 -12196 32708 -12188
rect 32716 -12196 32744 -12188
rect 32752 -12196 32772 -12188
rect 32808 -12188 32892 -12168
rect 32808 -12196 32828 -12188
rect 32836 -12196 32864 -12188
rect 32872 -12196 32892 -12188
rect 32928 -12188 33012 -12168
rect 32928 -12196 32948 -12188
rect 32956 -12196 32984 -12188
rect 32992 -12196 33012 -12188
rect 33048 -12188 33132 -12168
rect 33048 -12196 33068 -12188
rect 33076 -12196 33104 -12188
rect 33112 -12196 33132 -12188
rect 33168 -12188 33252 -12168
rect 33168 -12196 33188 -12188
rect 33196 -12196 33224 -12188
rect 33232 -12196 33252 -12188
rect 33288 -12188 33372 -12168
rect 33288 -12196 33308 -12188
rect 33316 -12196 33344 -12188
rect 33352 -12196 33372 -12188
rect 33408 -12188 33492 -12168
rect 33408 -12196 33428 -12188
rect 33436 -12196 33464 -12188
rect 33472 -12196 33492 -12188
rect 33528 -12188 33612 -12168
rect 33528 -12196 33548 -12188
rect 33556 -12196 33584 -12188
rect 33592 -12196 33612 -12188
rect 33648 -12188 33732 -12168
rect 33648 -12196 33668 -12188
rect 33676 -12196 33704 -12188
rect 33712 -12196 33732 -12188
rect 33768 -12188 33852 -12168
rect 33768 -12196 33788 -12188
rect 33796 -12196 33824 -12188
rect 33832 -12196 33852 -12188
rect 33888 -12188 33972 -12168
rect 33888 -12196 33908 -12188
rect 33916 -12196 33944 -12188
rect 33952 -12196 33972 -12188
rect 34008 -12188 34092 -12168
rect 34008 -12196 34028 -12188
rect 34036 -12196 34064 -12188
rect 34072 -12196 34092 -12188
rect 34128 -12188 34212 -12168
rect 34128 -12196 34148 -12188
rect 34156 -12196 34184 -12188
rect 34192 -12196 34212 -12188
rect 34248 -12188 34332 -12168
rect 34248 -12196 34268 -12188
rect 34276 -12196 34304 -12188
rect 34312 -12196 34332 -12188
rect 34368 -12188 34452 -12168
rect 34368 -12196 34388 -12188
rect 34396 -12196 34424 -12188
rect 34432 -12196 34452 -12188
rect 34488 -12188 34572 -12168
rect 34488 -12196 34508 -12188
rect 34516 -12196 34544 -12188
rect 34552 -12196 34572 -12188
rect 34608 -12188 34692 -12168
rect 34608 -12196 34628 -12188
rect 34636 -12196 34664 -12188
rect 34672 -12196 34692 -12188
rect 34728 -12188 34812 -12168
rect 34728 -12196 34748 -12188
rect 34756 -12196 34784 -12188
rect 34792 -12196 34812 -12188
rect 34848 -12188 34932 -12168
rect 34848 -12196 34868 -12188
rect 34876 -12196 34904 -12188
rect 34912 -12196 34932 -12188
rect 34968 -12188 35052 -12168
rect 34968 -12196 34988 -12188
rect 34996 -12196 35024 -12188
rect 35032 -12196 35052 -12188
rect 35088 -12188 35172 -12168
rect 35088 -12196 35108 -12188
rect 35116 -12196 35144 -12188
rect 35152 -12196 35172 -12188
rect 35208 -12188 35292 -12168
rect 35208 -12196 35228 -12188
rect 35236 -12196 35264 -12188
rect 35272 -12196 35292 -12188
rect 35328 -12188 35412 -12168
rect 35328 -12196 35348 -12188
rect 35356 -12196 35384 -12188
rect 35392 -12196 35412 -12188
rect 35448 -12188 35532 -12168
rect 35448 -12196 35468 -12188
rect 35476 -12196 35504 -12188
rect 35512 -12196 35532 -12188
rect 35568 -12188 35652 -12168
rect 35568 -12196 35588 -12188
rect 35596 -12196 35624 -12188
rect 35632 -12196 35652 -12188
rect 35688 -12188 35772 -12168
rect 35688 -12196 35708 -12188
rect 35716 -12196 35744 -12188
rect 35752 -12196 35772 -12188
rect 35808 -12188 35892 -12168
rect 35808 -12196 35828 -12188
rect 35836 -12196 35864 -12188
rect 35872 -12196 35892 -12188
rect 35928 -12188 36012 -12168
rect 35928 -12196 35948 -12188
rect 35956 -12196 35984 -12188
rect 35992 -12196 36012 -12188
rect 36048 -12188 36132 -12168
rect 36048 -12196 36068 -12188
rect 36076 -12196 36104 -12188
rect 36112 -12196 36132 -12188
rect 36168 -12188 36252 -12168
rect 36168 -12196 36188 -12188
rect 36196 -12196 36224 -12188
rect 36232 -12196 36252 -12188
rect 36288 -12188 36372 -12168
rect 36288 -12196 36308 -12188
rect 36316 -12196 36344 -12188
rect 36352 -12196 36372 -12188
rect 36408 -12188 36492 -12168
rect 36408 -12196 36428 -12188
rect 36436 -12196 36464 -12188
rect 36472 -12196 36492 -12188
rect 36528 -12188 36612 -12168
rect 36528 -12196 36548 -12188
rect 36556 -12196 36584 -12188
rect 36592 -12196 36612 -12188
rect 36648 -12188 36732 -12168
rect 36648 -12196 36668 -12188
rect 36676 -12196 36704 -12188
rect 36712 -12196 36732 -12188
rect 36768 -12188 36852 -12168
rect 36768 -12196 36788 -12188
rect 36796 -12196 36824 -12188
rect 36832 -12196 36852 -12188
rect 36888 -12188 36972 -12168
rect 36888 -12196 36908 -12188
rect 36916 -12196 36944 -12188
rect 36952 -12196 36972 -12188
rect 37008 -12188 37092 -12168
rect 37008 -12196 37028 -12188
rect 37036 -12196 37064 -12188
rect 37072 -12196 37092 -12188
rect 37128 -12188 37212 -12168
rect 37128 -12196 37148 -12188
rect 37156 -12196 37184 -12188
rect 37192 -12196 37212 -12188
rect 37248 -12188 37332 -12168
rect 37248 -12196 37268 -12188
rect 37276 -12196 37304 -12188
rect 37312 -12196 37332 -12188
rect 37368 -12188 37452 -12168
rect 37368 -12196 37388 -12188
rect 37396 -12196 37424 -12188
rect 37432 -12196 37452 -12188
rect 37488 -12188 37572 -12168
rect 37488 -12196 37508 -12188
rect 37516 -12196 37544 -12188
rect 37552 -12196 37572 -12188
rect 37608 -12188 37692 -12168
rect 37608 -12196 37628 -12188
rect 37636 -12196 37664 -12188
rect 37672 -12196 37692 -12188
rect 37728 -12188 37812 -12168
rect 37728 -12196 37748 -12188
rect 37756 -12196 37784 -12188
rect 37792 -12196 37812 -12188
rect 37848 -12188 37932 -12168
rect 37848 -12196 37868 -12188
rect 37876 -12196 37904 -12188
rect 37912 -12196 37932 -12188
rect 37968 -12188 38052 -12168
rect 37968 -12196 37988 -12188
rect 37996 -12196 38024 -12188
rect 38032 -12196 38052 -12188
rect 38088 -12188 38172 -12168
rect 38088 -12196 38108 -12188
rect 38116 -12196 38144 -12188
rect 38152 -12196 38172 -12188
rect 38208 -12188 38292 -12168
rect 38208 -12196 38228 -12188
rect 38236 -12196 38264 -12188
rect 38272 -12196 38292 -12188
rect 38328 -12188 38412 -12168
rect 38328 -12196 38348 -12188
rect 38356 -12196 38384 -12188
rect 38392 -12196 38412 -12188
rect 38448 -12188 38532 -12168
rect 38448 -12196 38468 -12188
rect 38476 -12196 38504 -12188
rect 38512 -12196 38532 -12188
rect 38568 -12188 38652 -12168
rect 38568 -12196 38588 -12188
rect 38596 -12196 38624 -12188
rect 38632 -12196 38652 -12188
rect 38688 -12188 38772 -12168
rect 38688 -12196 38708 -12188
rect 38716 -12196 38744 -12188
rect 38752 -12196 38772 -12188
rect 38808 -12188 38892 -12168
rect 38808 -12196 38828 -12188
rect 38836 -12196 38864 -12188
rect 38872 -12196 38892 -12188
rect 38928 -12188 39012 -12168
rect 38928 -12196 38948 -12188
rect 38956 -12196 38984 -12188
rect 38992 -12196 39012 -12188
rect 39048 -12188 39132 -12168
rect 39048 -12196 39068 -12188
rect 39076 -12196 39104 -12188
rect 39112 -12196 39132 -12188
rect 39168 -12188 39252 -12168
rect 39168 -12196 39188 -12188
rect 39196 -12196 39224 -12188
rect 39232 -12196 39252 -12188
rect 39288 -12188 39372 -12168
rect 39288 -12196 39308 -12188
rect 39316 -12196 39344 -12188
rect 39352 -12196 39372 -12188
rect 39408 -12188 39492 -12168
rect 39408 -12196 39428 -12188
rect 39436 -12196 39464 -12188
rect 39472 -12196 39492 -12188
rect 39528 -12188 39612 -12168
rect 39528 -12196 39548 -12188
rect 39556 -12196 39584 -12188
rect 39592 -12196 39612 -12188
rect 39648 -12188 39732 -12168
rect 39648 -12196 39668 -12188
rect 39676 -12196 39704 -12188
rect 39712 -12196 39732 -12188
rect 39768 -12188 39852 -12168
rect 39768 -12196 39788 -12188
rect 39796 -12196 39824 -12188
rect 39832 -12196 39852 -12188
rect 39888 -12188 39972 -12168
rect 39888 -12196 39908 -12188
rect 39916 -12196 39944 -12188
rect 39952 -12196 39972 -12188
rect 40008 -12188 40092 -12168
rect 40008 -12196 40028 -12188
rect 40036 -12196 40064 -12188
rect 40072 -12196 40092 -12188
rect 40128 -12188 40212 -12168
rect 40128 -12196 40148 -12188
rect 40156 -12196 40184 -12188
rect 40192 -12196 40212 -12188
rect 40248 -12188 40332 -12168
rect 40248 -12196 40268 -12188
rect 40276 -12196 40304 -12188
rect 40312 -12196 40332 -12188
rect 40368 -12188 40452 -12168
rect 40368 -12196 40388 -12188
rect 40396 -12196 40424 -12188
rect 40432 -12196 40452 -12188
rect 40488 -12188 40572 -12168
rect 40488 -12196 40508 -12188
rect 40516 -12196 40544 -12188
rect 40552 -12196 40572 -12188
rect 40608 -12188 40692 -12168
rect 40608 -12196 40628 -12188
rect 40636 -12196 40664 -12188
rect 40672 -12196 40692 -12188
rect 40728 -12188 40812 -12168
rect 40728 -12196 40748 -12188
rect 40756 -12196 40784 -12188
rect 40792 -12196 40812 -12188
rect 40848 -12188 40932 -12168
rect 40848 -12196 40868 -12188
rect 40876 -12196 40904 -12188
rect 40912 -12196 40932 -12188
rect 40968 -12188 41052 -12168
rect 40968 -12196 40988 -12188
rect 40996 -12196 41024 -12188
rect 41032 -12196 41052 -12188
rect 41088 -12188 41172 -12168
rect 41088 -12196 41108 -12188
rect 41116 -12196 41144 -12188
rect 41152 -12196 41172 -12188
rect 41208 -12188 41292 -12168
rect 41208 -12196 41228 -12188
rect 41236 -12196 41264 -12188
rect 41272 -12196 41292 -12188
rect 41328 -12188 41412 -12168
rect 41328 -12196 41348 -12188
rect 41356 -12196 41384 -12188
rect 41392 -12196 41412 -12188
rect 41448 -12188 41532 -12168
rect 41448 -12196 41468 -12188
rect 41476 -12196 41504 -12188
rect 41512 -12196 41532 -12188
rect 41568 -12188 41652 -12168
rect 41568 -12196 41588 -12188
rect 41596 -12196 41624 -12188
rect 41632 -12196 41652 -12188
rect 41688 -12188 41772 -12168
rect 41688 -12196 41708 -12188
rect 41716 -12196 41744 -12188
rect 41752 -12196 41772 -12188
rect 41808 -12188 41892 -12168
rect 41808 -12196 41828 -12188
rect 41836 -12196 41864 -12188
rect 41872 -12196 41892 -12188
rect 41928 -12188 42012 -12168
rect 41928 -12196 41948 -12188
rect 41956 -12196 41984 -12188
rect 41992 -12196 42012 -12188
rect 42048 -12188 42132 -12168
rect 42048 -12196 42068 -12188
rect 42076 -12196 42104 -12188
rect 42112 -12196 42132 -12188
rect 42168 -12188 42252 -12168
rect 42168 -12196 42188 -12188
rect 42196 -12196 42224 -12188
rect 42232 -12196 42252 -12188
rect 42288 -12188 42372 -12168
rect 42288 -12196 42308 -12188
rect 42316 -12196 42344 -12188
rect 42352 -12196 42372 -12188
rect 42408 -12188 42492 -12168
rect 42408 -12196 42428 -12188
rect 42436 -12196 42464 -12188
rect 42472 -12196 42492 -12188
rect 42528 -12188 42612 -12168
rect 42528 -12196 42548 -12188
rect 42556 -12196 42584 -12188
rect 42592 -12196 42612 -12188
rect 42648 -12188 42732 -12168
rect 42648 -12196 42668 -12188
rect 42676 -12196 42704 -12188
rect 42712 -12196 42732 -12188
rect 42768 -12188 42852 -12168
rect 42768 -12196 42788 -12188
rect 42796 -12196 42824 -12188
rect 42832 -12196 42852 -12188
rect 42888 -12188 42972 -12168
rect 42888 -12196 42908 -12188
rect 42916 -12196 42944 -12188
rect 42952 -12196 42972 -12188
rect 43008 -12188 43092 -12168
rect 43008 -12196 43028 -12188
rect 43036 -12196 43064 -12188
rect 43072 -12196 43092 -12188
rect 43128 -12188 43212 -12168
rect 43128 -12196 43148 -12188
rect 43156 -12196 43184 -12188
rect 43192 -12196 43212 -12188
rect 43248 -12188 43332 -12168
rect 43248 -12196 43268 -12188
rect 43276 -12196 43304 -12188
rect 43312 -12196 43332 -12188
rect 43368 -12188 43452 -12168
rect 43368 -12196 43388 -12188
rect 43396 -12196 43424 -12188
rect 43432 -12196 43452 -12188
rect 43488 -12188 43572 -12168
rect 43488 -12196 43508 -12188
rect 43516 -12196 43544 -12188
rect 43552 -12196 43572 -12188
rect 43608 -12188 43692 -12168
rect 43608 -12196 43628 -12188
rect 43636 -12196 43664 -12188
rect 43672 -12196 43692 -12188
rect 43728 -12188 43812 -12168
rect 43728 -12196 43748 -12188
rect 43756 -12196 43784 -12188
rect 43792 -12196 43812 -12188
rect 43848 -12188 43932 -12168
rect 43848 -12196 43868 -12188
rect 43876 -12196 43904 -12188
rect 43912 -12196 43932 -12188
rect 43968 -12188 44052 -12168
rect 43968 -12196 43988 -12188
rect 43996 -12196 44024 -12188
rect 44032 -12196 44052 -12188
rect 44088 -12188 44172 -12168
rect 44088 -12196 44108 -12188
rect 44116 -12196 44144 -12188
rect 44152 -12196 44172 -12188
rect 44208 -12188 44292 -12168
rect 44208 -12196 44228 -12188
rect 44236 -12196 44264 -12188
rect 44272 -12196 44292 -12188
rect 44328 -12188 44412 -12168
rect 44328 -12196 44348 -12188
rect 44356 -12196 44384 -12188
rect 44392 -12196 44412 -12188
rect 44448 -12188 44532 -12168
rect 44448 -12196 44468 -12188
rect 44476 -12196 44504 -12188
rect 44512 -12196 44532 -12188
rect 44568 -12188 44652 -12168
rect 44568 -12196 44588 -12188
rect 44596 -12196 44624 -12188
rect 44632 -12196 44652 -12188
rect 44688 -12188 44772 -12168
rect 44688 -12196 44708 -12188
rect 44716 -12196 44744 -12188
rect 44752 -12196 44772 -12188
rect 44808 -12188 44892 -12168
rect 44808 -12196 44828 -12188
rect 44836 -12196 44864 -12188
rect 44872 -12196 44892 -12188
rect 44928 -12188 45012 -12168
rect 44928 -12196 44948 -12188
rect 44956 -12196 44984 -12188
rect 44992 -12196 45012 -12188
rect 45048 -12188 45132 -12168
rect 45048 -12196 45068 -12188
rect 45076 -12196 45104 -12188
rect 45112 -12196 45132 -12188
rect 45168 -12188 45252 -12168
rect 45168 -12196 45188 -12188
rect 45196 -12196 45224 -12188
rect 45232 -12196 45252 -12188
rect 45288 -12188 45372 -12168
rect 45288 -12196 45308 -12188
rect 45316 -12196 45344 -12188
rect 45352 -12196 45372 -12188
rect 45408 -12188 45492 -12168
rect 45408 -12196 45428 -12188
rect 45436 -12196 45464 -12188
rect 45472 -12196 45492 -12188
rect 45528 -12188 45612 -12168
rect 45528 -12196 45548 -12188
rect 45556 -12196 45584 -12188
rect 45592 -12196 45612 -12188
rect 25876 -12224 25932 -12196
rect 25996 -12224 26052 -12196
rect 26116 -12224 26172 -12196
rect 26236 -12224 26292 -12196
rect 26356 -12224 26412 -12196
rect 26476 -12224 26532 -12196
rect 26596 -12224 26652 -12196
rect 26716 -12224 26772 -12196
rect 26836 -12224 26892 -12196
rect 26956 -12224 27012 -12196
rect 27076 -12224 27132 -12196
rect 27196 -12224 27252 -12196
rect 27316 -12224 27372 -12196
rect 27436 -12224 27492 -12196
rect 27556 -12224 27612 -12196
rect 27676 -12224 27732 -12196
rect 27796 -12224 27852 -12196
rect 27916 -12224 27972 -12196
rect 28036 -12224 28092 -12196
rect 28156 -12224 28212 -12196
rect 28276 -12224 28332 -12196
rect 28396 -12224 28452 -12196
rect 28516 -12224 28572 -12196
rect 28636 -12224 28692 -12196
rect 28756 -12224 28812 -12196
rect 28876 -12224 28932 -12196
rect 28996 -12224 29052 -12196
rect 29116 -12224 29172 -12196
rect 29236 -12224 29292 -12196
rect 29356 -12224 29412 -12196
rect 29476 -12224 29532 -12196
rect 29596 -12224 29652 -12196
rect 29716 -12224 29772 -12196
rect 29836 -12224 29892 -12196
rect 29956 -12224 30012 -12196
rect 30076 -12224 30132 -12196
rect 30196 -12224 30252 -12196
rect 30316 -12224 30372 -12196
rect 30436 -12224 30492 -12196
rect 30556 -12224 30612 -12196
rect 30676 -12224 30732 -12196
rect 30796 -12224 30852 -12196
rect 30916 -12224 30972 -12196
rect 31036 -12224 31092 -12196
rect 31156 -12224 31212 -12196
rect 31276 -12224 31332 -12196
rect 31396 -12224 31452 -12196
rect 31516 -12224 31572 -12196
rect 31636 -12224 31692 -12196
rect 31756 -12224 31812 -12196
rect 31876 -12224 31932 -12196
rect 31996 -12224 32052 -12196
rect 32116 -12224 32172 -12196
rect 32236 -12224 32292 -12196
rect 32356 -12224 32412 -12196
rect 32476 -12224 32532 -12196
rect 32596 -12224 32652 -12196
rect 32716 -12224 32772 -12196
rect 32836 -12224 32892 -12196
rect 32956 -12224 33012 -12196
rect 33076 -12224 33132 -12196
rect 33196 -12224 33252 -12196
rect 33316 -12224 33372 -12196
rect 33436 -12224 33492 -12196
rect 33556 -12224 33612 -12196
rect 33676 -12224 33732 -12196
rect 33796 -12224 33852 -12196
rect 33916 -12224 33972 -12196
rect 34036 -12224 34092 -12196
rect 34156 -12224 34212 -12196
rect 34276 -12224 34332 -12196
rect 34396 -12224 34452 -12196
rect 34516 -12224 34572 -12196
rect 34636 -12224 34692 -12196
rect 34756 -12224 34812 -12196
rect 34876 -12224 34932 -12196
rect 34996 -12224 35052 -12196
rect 35116 -12224 35172 -12196
rect 35236 -12224 35292 -12196
rect 35356 -12224 35412 -12196
rect 35476 -12224 35532 -12196
rect 35596 -12224 35652 -12196
rect 35716 -12224 35772 -12196
rect 35836 -12224 35892 -12196
rect 35956 -12224 36012 -12196
rect 36076 -12224 36132 -12196
rect 36196 -12224 36252 -12196
rect 36316 -12224 36372 -12196
rect 36436 -12224 36492 -12196
rect 36556 -12224 36612 -12196
rect 36676 -12224 36732 -12196
rect 36796 -12224 36852 -12196
rect 36916 -12224 36972 -12196
rect 37036 -12224 37092 -12196
rect 37156 -12224 37212 -12196
rect 37276 -12224 37332 -12196
rect 37396 -12224 37452 -12196
rect 37516 -12224 37572 -12196
rect 37636 -12224 37692 -12196
rect 37756 -12224 37812 -12196
rect 37876 -12224 37932 -12196
rect 37996 -12224 38052 -12196
rect 38116 -12224 38172 -12196
rect 38236 -12224 38292 -12196
rect 38356 -12224 38412 -12196
rect 38476 -12224 38532 -12196
rect 38596 -12224 38652 -12196
rect 38716 -12224 38772 -12196
rect 38836 -12224 38892 -12196
rect 38956 -12224 39012 -12196
rect 39076 -12224 39132 -12196
rect 39196 -12224 39252 -12196
rect 39316 -12224 39372 -12196
rect 39436 -12224 39492 -12196
rect 39556 -12224 39612 -12196
rect 39676 -12224 39732 -12196
rect 39796 -12224 39852 -12196
rect 39916 -12224 39972 -12196
rect 40036 -12224 40092 -12196
rect 40156 -12224 40212 -12196
rect 40276 -12224 40332 -12196
rect 40396 -12224 40452 -12196
rect 40516 -12224 40572 -12196
rect 40636 -12224 40692 -12196
rect 40756 -12224 40812 -12196
rect 40876 -12224 40932 -12196
rect 40996 -12224 41052 -12196
rect 41116 -12224 41172 -12196
rect 41236 -12224 41292 -12196
rect 41356 -12224 41412 -12196
rect 41476 -12224 41532 -12196
rect 41596 -12224 41652 -12196
rect 41716 -12224 41772 -12196
rect 41836 -12224 41892 -12196
rect 41956 -12224 42012 -12196
rect 42076 -12224 42132 -12196
rect 42196 -12224 42252 -12196
rect 42316 -12224 42372 -12196
rect 42436 -12224 42492 -12196
rect 42556 -12224 42612 -12196
rect 42676 -12224 42732 -12196
rect 42796 -12224 42852 -12196
rect 42916 -12224 42972 -12196
rect 43036 -12224 43092 -12196
rect 43156 -12224 43212 -12196
rect 43276 -12224 43332 -12196
rect 43396 -12224 43452 -12196
rect 43516 -12224 43572 -12196
rect 43636 -12224 43692 -12196
rect 43756 -12224 43812 -12196
rect 43876 -12224 43932 -12196
rect 43996 -12224 44052 -12196
rect 44116 -12224 44172 -12196
rect 44236 -12224 44292 -12196
rect 44356 -12224 44412 -12196
rect 44476 -12224 44532 -12196
rect 44596 -12224 44652 -12196
rect 44716 -12224 44772 -12196
rect 44836 -12224 44892 -12196
rect 44956 -12224 45012 -12196
rect 45076 -12224 45132 -12196
rect 45196 -12224 45252 -12196
rect 45316 -12224 45372 -12196
rect 45436 -12224 45492 -12196
rect 45556 -12224 45612 -12196
rect 25848 -12368 25932 -12348
rect 25848 -12376 25868 -12368
rect 25876 -12376 25904 -12368
rect 25912 -12376 25932 -12368
rect 25968 -12368 26052 -12348
rect 25968 -12376 25988 -12368
rect 25996 -12376 26024 -12368
rect 26032 -12376 26052 -12368
rect 26088 -12368 26172 -12348
rect 26088 -12376 26108 -12368
rect 26116 -12376 26144 -12368
rect 26152 -12376 26172 -12368
rect 26208 -12368 26292 -12348
rect 26208 -12376 26228 -12368
rect 26236 -12376 26264 -12368
rect 26272 -12376 26292 -12368
rect 26328 -12368 26412 -12348
rect 26328 -12376 26348 -12368
rect 26356 -12376 26384 -12368
rect 26392 -12376 26412 -12368
rect 26448 -12368 26532 -12348
rect 26448 -12376 26468 -12368
rect 26476 -12376 26504 -12368
rect 26512 -12376 26532 -12368
rect 26568 -12368 26652 -12348
rect 26568 -12376 26588 -12368
rect 26596 -12376 26624 -12368
rect 26632 -12376 26652 -12368
rect 26688 -12368 26772 -12348
rect 26688 -12376 26708 -12368
rect 26716 -12376 26744 -12368
rect 26752 -12376 26772 -12368
rect 26808 -12368 26892 -12348
rect 26808 -12376 26828 -12368
rect 26836 -12376 26864 -12368
rect 26872 -12376 26892 -12368
rect 26928 -12368 27012 -12348
rect 26928 -12376 26948 -12368
rect 26956 -12376 26984 -12368
rect 26992 -12376 27012 -12368
rect 27048 -12368 27132 -12348
rect 27048 -12376 27068 -12368
rect 27076 -12376 27104 -12368
rect 27112 -12376 27132 -12368
rect 27168 -12368 27252 -12348
rect 27168 -12376 27188 -12368
rect 27196 -12376 27224 -12368
rect 27232 -12376 27252 -12368
rect 27288 -12368 27372 -12348
rect 27288 -12376 27308 -12368
rect 27316 -12376 27344 -12368
rect 27352 -12376 27372 -12368
rect 27408 -12368 27492 -12348
rect 27408 -12376 27428 -12368
rect 27436 -12376 27464 -12368
rect 27472 -12376 27492 -12368
rect 27528 -12368 27612 -12348
rect 27528 -12376 27548 -12368
rect 27556 -12376 27584 -12368
rect 27592 -12376 27612 -12368
rect 27648 -12368 27732 -12348
rect 27648 -12376 27668 -12368
rect 27676 -12376 27704 -12368
rect 27712 -12376 27732 -12368
rect 27768 -12368 27852 -12348
rect 27768 -12376 27788 -12368
rect 27796 -12376 27824 -12368
rect 27832 -12376 27852 -12368
rect 27888 -12368 27972 -12348
rect 27888 -12376 27908 -12368
rect 27916 -12376 27944 -12368
rect 27952 -12376 27972 -12368
rect 28008 -12368 28092 -12348
rect 28008 -12376 28028 -12368
rect 28036 -12376 28064 -12368
rect 28072 -12376 28092 -12368
rect 28128 -12368 28212 -12348
rect 28128 -12376 28148 -12368
rect 28156 -12376 28184 -12368
rect 28192 -12376 28212 -12368
rect 28248 -12368 28332 -12348
rect 28248 -12376 28268 -12368
rect 28276 -12376 28304 -12368
rect 28312 -12376 28332 -12368
rect 28368 -12368 28452 -12348
rect 28368 -12376 28388 -12368
rect 28396 -12376 28424 -12368
rect 28432 -12376 28452 -12368
rect 28488 -12368 28572 -12348
rect 28488 -12376 28508 -12368
rect 28516 -12376 28544 -12368
rect 28552 -12376 28572 -12368
rect 28608 -12368 28692 -12348
rect 28608 -12376 28628 -12368
rect 28636 -12376 28664 -12368
rect 28672 -12376 28692 -12368
rect 28728 -12368 28812 -12348
rect 28728 -12376 28748 -12368
rect 28756 -12376 28784 -12368
rect 28792 -12376 28812 -12368
rect 28848 -12368 28932 -12348
rect 28848 -12376 28868 -12368
rect 28876 -12376 28904 -12368
rect 28912 -12376 28932 -12368
rect 28968 -12368 29052 -12348
rect 28968 -12376 28988 -12368
rect 28996 -12376 29024 -12368
rect 29032 -12376 29052 -12368
rect 29088 -12368 29172 -12348
rect 29088 -12376 29108 -12368
rect 29116 -12376 29144 -12368
rect 29152 -12376 29172 -12368
rect 29208 -12368 29292 -12348
rect 29208 -12376 29228 -12368
rect 29236 -12376 29264 -12368
rect 29272 -12376 29292 -12368
rect 29328 -12368 29412 -12348
rect 29328 -12376 29348 -12368
rect 29356 -12376 29384 -12368
rect 29392 -12376 29412 -12368
rect 29448 -12368 29532 -12348
rect 29448 -12376 29468 -12368
rect 29476 -12376 29504 -12368
rect 29512 -12376 29532 -12368
rect 29568 -12368 29652 -12348
rect 29568 -12376 29588 -12368
rect 29596 -12376 29624 -12368
rect 29632 -12376 29652 -12368
rect 29688 -12368 29772 -12348
rect 29688 -12376 29708 -12368
rect 29716 -12376 29744 -12368
rect 29752 -12376 29772 -12368
rect 29808 -12368 29892 -12348
rect 29808 -12376 29828 -12368
rect 29836 -12376 29864 -12368
rect 29872 -12376 29892 -12368
rect 29928 -12368 30012 -12348
rect 29928 -12376 29948 -12368
rect 29956 -12376 29984 -12368
rect 29992 -12376 30012 -12368
rect 30048 -12368 30132 -12348
rect 30048 -12376 30068 -12368
rect 30076 -12376 30104 -12368
rect 30112 -12376 30132 -12368
rect 30168 -12368 30252 -12348
rect 30168 -12376 30188 -12368
rect 30196 -12376 30224 -12368
rect 30232 -12376 30252 -12368
rect 30288 -12368 30372 -12348
rect 30288 -12376 30308 -12368
rect 30316 -12376 30344 -12368
rect 30352 -12376 30372 -12368
rect 30408 -12368 30492 -12348
rect 30408 -12376 30428 -12368
rect 30436 -12376 30464 -12368
rect 30472 -12376 30492 -12368
rect 30528 -12368 30612 -12348
rect 30528 -12376 30548 -12368
rect 30556 -12376 30584 -12368
rect 30592 -12376 30612 -12368
rect 30648 -12368 30732 -12348
rect 30648 -12376 30668 -12368
rect 30676 -12376 30704 -12368
rect 30712 -12376 30732 -12368
rect 30768 -12368 30852 -12348
rect 30768 -12376 30788 -12368
rect 30796 -12376 30824 -12368
rect 30832 -12376 30852 -12368
rect 30888 -12368 30972 -12348
rect 30888 -12376 30908 -12368
rect 30916 -12376 30944 -12368
rect 30952 -12376 30972 -12368
rect 31008 -12368 31092 -12348
rect 31008 -12376 31028 -12368
rect 31036 -12376 31064 -12368
rect 31072 -12376 31092 -12368
rect 31128 -12368 31212 -12348
rect 31128 -12376 31148 -12368
rect 31156 -12376 31184 -12368
rect 31192 -12376 31212 -12368
rect 31248 -12368 31332 -12348
rect 31248 -12376 31268 -12368
rect 31276 -12376 31304 -12368
rect 31312 -12376 31332 -12368
rect 31368 -12368 31452 -12348
rect 31368 -12376 31388 -12368
rect 31396 -12376 31424 -12368
rect 31432 -12376 31452 -12368
rect 31488 -12368 31572 -12348
rect 31488 -12376 31508 -12368
rect 31516 -12376 31544 -12368
rect 31552 -12376 31572 -12368
rect 31608 -12368 31692 -12348
rect 31608 -12376 31628 -12368
rect 31636 -12376 31664 -12368
rect 31672 -12376 31692 -12368
rect 31728 -12368 31812 -12348
rect 31728 -12376 31748 -12368
rect 31756 -12376 31784 -12368
rect 31792 -12376 31812 -12368
rect 31848 -12368 31932 -12348
rect 31848 -12376 31868 -12368
rect 31876 -12376 31904 -12368
rect 31912 -12376 31932 -12368
rect 31968 -12368 32052 -12348
rect 31968 -12376 31988 -12368
rect 31996 -12376 32024 -12368
rect 32032 -12376 32052 -12368
rect 32088 -12368 32172 -12348
rect 32088 -12376 32108 -12368
rect 32116 -12376 32144 -12368
rect 32152 -12376 32172 -12368
rect 32208 -12368 32292 -12348
rect 32208 -12376 32228 -12368
rect 32236 -12376 32264 -12368
rect 32272 -12376 32292 -12368
rect 32328 -12368 32412 -12348
rect 32328 -12376 32348 -12368
rect 32356 -12376 32384 -12368
rect 32392 -12376 32412 -12368
rect 32448 -12368 32532 -12348
rect 32448 -12376 32468 -12368
rect 32476 -12376 32504 -12368
rect 32512 -12376 32532 -12368
rect 32568 -12368 32652 -12348
rect 32568 -12376 32588 -12368
rect 32596 -12376 32624 -12368
rect 32632 -12376 32652 -12368
rect 32688 -12368 32772 -12348
rect 32688 -12376 32708 -12368
rect 32716 -12376 32744 -12368
rect 32752 -12376 32772 -12368
rect 32808 -12368 32892 -12348
rect 32808 -12376 32828 -12368
rect 32836 -12376 32864 -12368
rect 32872 -12376 32892 -12368
rect 32928 -12368 33012 -12348
rect 32928 -12376 32948 -12368
rect 32956 -12376 32984 -12368
rect 32992 -12376 33012 -12368
rect 33048 -12368 33132 -12348
rect 33048 -12376 33068 -12368
rect 33076 -12376 33104 -12368
rect 33112 -12376 33132 -12368
rect 33168 -12368 33252 -12348
rect 33168 -12376 33188 -12368
rect 33196 -12376 33224 -12368
rect 33232 -12376 33252 -12368
rect 33288 -12368 33372 -12348
rect 33288 -12376 33308 -12368
rect 33316 -12376 33344 -12368
rect 33352 -12376 33372 -12368
rect 33408 -12368 33492 -12348
rect 33408 -12376 33428 -12368
rect 33436 -12376 33464 -12368
rect 33472 -12376 33492 -12368
rect 33528 -12368 33612 -12348
rect 33528 -12376 33548 -12368
rect 33556 -12376 33584 -12368
rect 33592 -12376 33612 -12368
rect 33648 -12368 33732 -12348
rect 33648 -12376 33668 -12368
rect 33676 -12376 33704 -12368
rect 33712 -12376 33732 -12368
rect 33768 -12368 33852 -12348
rect 33768 -12376 33788 -12368
rect 33796 -12376 33824 -12368
rect 33832 -12376 33852 -12368
rect 33888 -12368 33972 -12348
rect 33888 -12376 33908 -12368
rect 33916 -12376 33944 -12368
rect 33952 -12376 33972 -12368
rect 34008 -12368 34092 -12348
rect 34008 -12376 34028 -12368
rect 34036 -12376 34064 -12368
rect 34072 -12376 34092 -12368
rect 34128 -12368 34212 -12348
rect 34128 -12376 34148 -12368
rect 34156 -12376 34184 -12368
rect 34192 -12376 34212 -12368
rect 34248 -12368 34332 -12348
rect 34248 -12376 34268 -12368
rect 34276 -12376 34304 -12368
rect 34312 -12376 34332 -12368
rect 34368 -12368 34452 -12348
rect 34368 -12376 34388 -12368
rect 34396 -12376 34424 -12368
rect 34432 -12376 34452 -12368
rect 34488 -12368 34572 -12348
rect 34488 -12376 34508 -12368
rect 34516 -12376 34544 -12368
rect 34552 -12376 34572 -12368
rect 34608 -12368 34692 -12348
rect 34608 -12376 34628 -12368
rect 34636 -12376 34664 -12368
rect 34672 -12376 34692 -12368
rect 34728 -12368 34812 -12348
rect 34728 -12376 34748 -12368
rect 34756 -12376 34784 -12368
rect 34792 -12376 34812 -12368
rect 34848 -12368 34932 -12348
rect 34848 -12376 34868 -12368
rect 34876 -12376 34904 -12368
rect 34912 -12376 34932 -12368
rect 34968 -12368 35052 -12348
rect 34968 -12376 34988 -12368
rect 34996 -12376 35024 -12368
rect 35032 -12376 35052 -12368
rect 35088 -12368 35172 -12348
rect 35088 -12376 35108 -12368
rect 35116 -12376 35144 -12368
rect 35152 -12376 35172 -12368
rect 35208 -12368 35292 -12348
rect 35208 -12376 35228 -12368
rect 35236 -12376 35264 -12368
rect 35272 -12376 35292 -12368
rect 35328 -12368 35412 -12348
rect 35328 -12376 35348 -12368
rect 35356 -12376 35384 -12368
rect 35392 -12376 35412 -12368
rect 35448 -12368 35532 -12348
rect 35448 -12376 35468 -12368
rect 35476 -12376 35504 -12368
rect 35512 -12376 35532 -12368
rect 35568 -12368 35652 -12348
rect 35568 -12376 35588 -12368
rect 35596 -12376 35624 -12368
rect 35632 -12376 35652 -12368
rect 35688 -12368 35772 -12348
rect 35688 -12376 35708 -12368
rect 35716 -12376 35744 -12368
rect 35752 -12376 35772 -12368
rect 35808 -12368 35892 -12348
rect 35808 -12376 35828 -12368
rect 35836 -12376 35864 -12368
rect 35872 -12376 35892 -12368
rect 35928 -12368 36012 -12348
rect 35928 -12376 35948 -12368
rect 35956 -12376 35984 -12368
rect 35992 -12376 36012 -12368
rect 36048 -12368 36132 -12348
rect 36048 -12376 36068 -12368
rect 36076 -12376 36104 -12368
rect 36112 -12376 36132 -12368
rect 36168 -12368 36252 -12348
rect 36168 -12376 36188 -12368
rect 36196 -12376 36224 -12368
rect 36232 -12376 36252 -12368
rect 36288 -12368 36372 -12348
rect 36288 -12376 36308 -12368
rect 36316 -12376 36344 -12368
rect 36352 -12376 36372 -12368
rect 36408 -12368 36492 -12348
rect 36408 -12376 36428 -12368
rect 36436 -12376 36464 -12368
rect 36472 -12376 36492 -12368
rect 36528 -12368 36612 -12348
rect 36528 -12376 36548 -12368
rect 36556 -12376 36584 -12368
rect 36592 -12376 36612 -12368
rect 36648 -12368 36732 -12348
rect 36648 -12376 36668 -12368
rect 36676 -12376 36704 -12368
rect 36712 -12376 36732 -12368
rect 36768 -12368 36852 -12348
rect 36768 -12376 36788 -12368
rect 36796 -12376 36824 -12368
rect 36832 -12376 36852 -12368
rect 36888 -12368 36972 -12348
rect 36888 -12376 36908 -12368
rect 36916 -12376 36944 -12368
rect 36952 -12376 36972 -12368
rect 37008 -12368 37092 -12348
rect 37008 -12376 37028 -12368
rect 37036 -12376 37064 -12368
rect 37072 -12376 37092 -12368
rect 37128 -12368 37212 -12348
rect 37128 -12376 37148 -12368
rect 37156 -12376 37184 -12368
rect 37192 -12376 37212 -12368
rect 37248 -12368 37332 -12348
rect 37248 -12376 37268 -12368
rect 37276 -12376 37304 -12368
rect 37312 -12376 37332 -12368
rect 37368 -12368 37452 -12348
rect 37368 -12376 37388 -12368
rect 37396 -12376 37424 -12368
rect 37432 -12376 37452 -12368
rect 37488 -12368 37572 -12348
rect 37488 -12376 37508 -12368
rect 37516 -12376 37544 -12368
rect 37552 -12376 37572 -12368
rect 37608 -12368 37692 -12348
rect 37608 -12376 37628 -12368
rect 37636 -12376 37664 -12368
rect 37672 -12376 37692 -12368
rect 37728 -12368 37812 -12348
rect 37728 -12376 37748 -12368
rect 37756 -12376 37784 -12368
rect 37792 -12376 37812 -12368
rect 37848 -12368 37932 -12348
rect 37848 -12376 37868 -12368
rect 37876 -12376 37904 -12368
rect 37912 -12376 37932 -12368
rect 37968 -12368 38052 -12348
rect 37968 -12376 37988 -12368
rect 37996 -12376 38024 -12368
rect 38032 -12376 38052 -12368
rect 38088 -12368 38172 -12348
rect 38088 -12376 38108 -12368
rect 38116 -12376 38144 -12368
rect 38152 -12376 38172 -12368
rect 38208 -12368 38292 -12348
rect 38208 -12376 38228 -12368
rect 38236 -12376 38264 -12368
rect 38272 -12376 38292 -12368
rect 38328 -12368 38412 -12348
rect 38328 -12376 38348 -12368
rect 38356 -12376 38384 -12368
rect 38392 -12376 38412 -12368
rect 38448 -12368 38532 -12348
rect 38448 -12376 38468 -12368
rect 38476 -12376 38504 -12368
rect 38512 -12376 38532 -12368
rect 38568 -12368 38652 -12348
rect 38568 -12376 38588 -12368
rect 38596 -12376 38624 -12368
rect 38632 -12376 38652 -12368
rect 38688 -12368 38772 -12348
rect 38688 -12376 38708 -12368
rect 38716 -12376 38744 -12368
rect 38752 -12376 38772 -12368
rect 38808 -12368 38892 -12348
rect 38808 -12376 38828 -12368
rect 38836 -12376 38864 -12368
rect 38872 -12376 38892 -12368
rect 38928 -12368 39012 -12348
rect 38928 -12376 38948 -12368
rect 38956 -12376 38984 -12368
rect 38992 -12376 39012 -12368
rect 39048 -12368 39132 -12348
rect 39048 -12376 39068 -12368
rect 39076 -12376 39104 -12368
rect 39112 -12376 39132 -12368
rect 39168 -12368 39252 -12348
rect 39168 -12376 39188 -12368
rect 39196 -12376 39224 -12368
rect 39232 -12376 39252 -12368
rect 39288 -12368 39372 -12348
rect 39288 -12376 39308 -12368
rect 39316 -12376 39344 -12368
rect 39352 -12376 39372 -12368
rect 39408 -12368 39492 -12348
rect 39408 -12376 39428 -12368
rect 39436 -12376 39464 -12368
rect 39472 -12376 39492 -12368
rect 39528 -12368 39612 -12348
rect 39528 -12376 39548 -12368
rect 39556 -12376 39584 -12368
rect 39592 -12376 39612 -12368
rect 39648 -12368 39732 -12348
rect 39648 -12376 39668 -12368
rect 39676 -12376 39704 -12368
rect 39712 -12376 39732 -12368
rect 39768 -12368 39852 -12348
rect 39768 -12376 39788 -12368
rect 39796 -12376 39824 -12368
rect 39832 -12376 39852 -12368
rect 39888 -12368 39972 -12348
rect 39888 -12376 39908 -12368
rect 39916 -12376 39944 -12368
rect 39952 -12376 39972 -12368
rect 40008 -12368 40092 -12348
rect 40008 -12376 40028 -12368
rect 40036 -12376 40064 -12368
rect 40072 -12376 40092 -12368
rect 40128 -12368 40212 -12348
rect 40128 -12376 40148 -12368
rect 40156 -12376 40184 -12368
rect 40192 -12376 40212 -12368
rect 40248 -12368 40332 -12348
rect 40248 -12376 40268 -12368
rect 40276 -12376 40304 -12368
rect 40312 -12376 40332 -12368
rect 40368 -12368 40452 -12348
rect 40368 -12376 40388 -12368
rect 40396 -12376 40424 -12368
rect 40432 -12376 40452 -12368
rect 40488 -12368 40572 -12348
rect 40488 -12376 40508 -12368
rect 40516 -12376 40544 -12368
rect 40552 -12376 40572 -12368
rect 40608 -12368 40692 -12348
rect 40608 -12376 40628 -12368
rect 40636 -12376 40664 -12368
rect 40672 -12376 40692 -12368
rect 40728 -12368 40812 -12348
rect 40728 -12376 40748 -12368
rect 40756 -12376 40784 -12368
rect 40792 -12376 40812 -12368
rect 40848 -12368 40932 -12348
rect 40848 -12376 40868 -12368
rect 40876 -12376 40904 -12368
rect 40912 -12376 40932 -12368
rect 40968 -12368 41052 -12348
rect 40968 -12376 40988 -12368
rect 40996 -12376 41024 -12368
rect 41032 -12376 41052 -12368
rect 41088 -12368 41172 -12348
rect 41088 -12376 41108 -12368
rect 41116 -12376 41144 -12368
rect 41152 -12376 41172 -12368
rect 41208 -12368 41292 -12348
rect 41208 -12376 41228 -12368
rect 41236 -12376 41264 -12368
rect 41272 -12376 41292 -12368
rect 41328 -12368 41412 -12348
rect 41328 -12376 41348 -12368
rect 41356 -12376 41384 -12368
rect 41392 -12376 41412 -12368
rect 41448 -12368 41532 -12348
rect 41448 -12376 41468 -12368
rect 41476 -12376 41504 -12368
rect 41512 -12376 41532 -12368
rect 41568 -12368 41652 -12348
rect 41568 -12376 41588 -12368
rect 41596 -12376 41624 -12368
rect 41632 -12376 41652 -12368
rect 41688 -12368 41772 -12348
rect 41688 -12376 41708 -12368
rect 41716 -12376 41744 -12368
rect 41752 -12376 41772 -12368
rect 41808 -12368 41892 -12348
rect 41808 -12376 41828 -12368
rect 41836 -12376 41864 -12368
rect 41872 -12376 41892 -12368
rect 41928 -12368 42012 -12348
rect 41928 -12376 41948 -12368
rect 41956 -12376 41984 -12368
rect 41992 -12376 42012 -12368
rect 42048 -12368 42132 -12348
rect 42048 -12376 42068 -12368
rect 42076 -12376 42104 -12368
rect 42112 -12376 42132 -12368
rect 42168 -12368 42252 -12348
rect 42168 -12376 42188 -12368
rect 42196 -12376 42224 -12368
rect 42232 -12376 42252 -12368
rect 42288 -12368 42372 -12348
rect 42288 -12376 42308 -12368
rect 42316 -12376 42344 -12368
rect 42352 -12376 42372 -12368
rect 42408 -12368 42492 -12348
rect 42408 -12376 42428 -12368
rect 42436 -12376 42464 -12368
rect 42472 -12376 42492 -12368
rect 42528 -12368 42612 -12348
rect 42528 -12376 42548 -12368
rect 42556 -12376 42584 -12368
rect 42592 -12376 42612 -12368
rect 42648 -12368 42732 -12348
rect 42648 -12376 42668 -12368
rect 42676 -12376 42704 -12368
rect 42712 -12376 42732 -12368
rect 42768 -12368 42852 -12348
rect 42768 -12376 42788 -12368
rect 42796 -12376 42824 -12368
rect 42832 -12376 42852 -12368
rect 42888 -12368 42972 -12348
rect 42888 -12376 42908 -12368
rect 42916 -12376 42944 -12368
rect 42952 -12376 42972 -12368
rect 43008 -12368 43092 -12348
rect 43008 -12376 43028 -12368
rect 43036 -12376 43064 -12368
rect 43072 -12376 43092 -12368
rect 43128 -12368 43212 -12348
rect 43128 -12376 43148 -12368
rect 43156 -12376 43184 -12368
rect 43192 -12376 43212 -12368
rect 43248 -12368 43332 -12348
rect 43248 -12376 43268 -12368
rect 43276 -12376 43304 -12368
rect 43312 -12376 43332 -12368
rect 43368 -12368 43452 -12348
rect 43368 -12376 43388 -12368
rect 43396 -12376 43424 -12368
rect 43432 -12376 43452 -12368
rect 43488 -12368 43572 -12348
rect 43488 -12376 43508 -12368
rect 43516 -12376 43544 -12368
rect 43552 -12376 43572 -12368
rect 43608 -12368 43692 -12348
rect 43608 -12376 43628 -12368
rect 43636 -12376 43664 -12368
rect 43672 -12376 43692 -12368
rect 43728 -12368 43812 -12348
rect 43728 -12376 43748 -12368
rect 43756 -12376 43784 -12368
rect 43792 -12376 43812 -12368
rect 43848 -12368 43932 -12348
rect 43848 -12376 43868 -12368
rect 43876 -12376 43904 -12368
rect 43912 -12376 43932 -12368
rect 43968 -12368 44052 -12348
rect 43968 -12376 43988 -12368
rect 43996 -12376 44024 -12368
rect 44032 -12376 44052 -12368
rect 44088 -12368 44172 -12348
rect 44088 -12376 44108 -12368
rect 44116 -12376 44144 -12368
rect 44152 -12376 44172 -12368
rect 44208 -12368 44292 -12348
rect 44208 -12376 44228 -12368
rect 44236 -12376 44264 -12368
rect 44272 -12376 44292 -12368
rect 44328 -12368 44412 -12348
rect 44328 -12376 44348 -12368
rect 44356 -12376 44384 -12368
rect 44392 -12376 44412 -12368
rect 44448 -12368 44532 -12348
rect 44448 -12376 44468 -12368
rect 44476 -12376 44504 -12368
rect 44512 -12376 44532 -12368
rect 44568 -12368 44652 -12348
rect 44568 -12376 44588 -12368
rect 44596 -12376 44624 -12368
rect 44632 -12376 44652 -12368
rect 44688 -12368 44772 -12348
rect 44688 -12376 44708 -12368
rect 44716 -12376 44744 -12368
rect 44752 -12376 44772 -12368
rect 44808 -12368 44892 -12348
rect 44808 -12376 44828 -12368
rect 44836 -12376 44864 -12368
rect 44872 -12376 44892 -12368
rect 44928 -12368 45012 -12348
rect 44928 -12376 44948 -12368
rect 44956 -12376 44984 -12368
rect 44992 -12376 45012 -12368
rect 45048 -12368 45132 -12348
rect 45048 -12376 45068 -12368
rect 45076 -12376 45104 -12368
rect 45112 -12376 45132 -12368
rect 45168 -12368 45252 -12348
rect 45168 -12376 45188 -12368
rect 45196 -12376 45224 -12368
rect 45232 -12376 45252 -12368
rect 45288 -12368 45372 -12348
rect 45288 -12376 45308 -12368
rect 45316 -12376 45344 -12368
rect 45352 -12376 45372 -12368
rect 45408 -12368 45492 -12348
rect 45408 -12376 45428 -12368
rect 45436 -12376 45464 -12368
rect 45472 -12376 45492 -12368
rect 45528 -12368 45612 -12348
rect 45528 -12376 45548 -12368
rect 45556 -12376 45584 -12368
rect 45592 -12376 45612 -12368
rect 25876 -12404 25932 -12376
rect 25996 -12404 26052 -12376
rect 26116 -12404 26172 -12376
rect 26236 -12404 26292 -12376
rect 26356 -12404 26412 -12376
rect 26476 -12404 26532 -12376
rect 26596 -12404 26652 -12376
rect 26716 -12404 26772 -12376
rect 26836 -12404 26892 -12376
rect 26956 -12404 27012 -12376
rect 27076 -12404 27132 -12376
rect 27196 -12404 27252 -12376
rect 27316 -12404 27372 -12376
rect 27436 -12404 27492 -12376
rect 27556 -12404 27612 -12376
rect 27676 -12404 27732 -12376
rect 27796 -12404 27852 -12376
rect 27916 -12404 27972 -12376
rect 28036 -12404 28092 -12376
rect 28156 -12404 28212 -12376
rect 28276 -12404 28332 -12376
rect 28396 -12404 28452 -12376
rect 28516 -12404 28572 -12376
rect 28636 -12404 28692 -12376
rect 28756 -12404 28812 -12376
rect 28876 -12404 28932 -12376
rect 28996 -12404 29052 -12376
rect 29116 -12404 29172 -12376
rect 29236 -12404 29292 -12376
rect 29356 -12404 29412 -12376
rect 29476 -12404 29532 -12376
rect 29596 -12404 29652 -12376
rect 29716 -12404 29772 -12376
rect 29836 -12404 29892 -12376
rect 29956 -12404 30012 -12376
rect 30076 -12404 30132 -12376
rect 30196 -12404 30252 -12376
rect 30316 -12404 30372 -12376
rect 30436 -12404 30492 -12376
rect 30556 -12404 30612 -12376
rect 30676 -12404 30732 -12376
rect 30796 -12404 30852 -12376
rect 30916 -12404 30972 -12376
rect 31036 -12404 31092 -12376
rect 31156 -12404 31212 -12376
rect 31276 -12404 31332 -12376
rect 31396 -12404 31452 -12376
rect 31516 -12404 31572 -12376
rect 31636 -12404 31692 -12376
rect 31756 -12404 31812 -12376
rect 31876 -12404 31932 -12376
rect 31996 -12404 32052 -12376
rect 32116 -12404 32172 -12376
rect 32236 -12404 32292 -12376
rect 32356 -12404 32412 -12376
rect 32476 -12404 32532 -12376
rect 32596 -12404 32652 -12376
rect 32716 -12404 32772 -12376
rect 32836 -12404 32892 -12376
rect 32956 -12404 33012 -12376
rect 33076 -12404 33132 -12376
rect 33196 -12404 33252 -12376
rect 33316 -12404 33372 -12376
rect 33436 -12404 33492 -12376
rect 33556 -12404 33612 -12376
rect 33676 -12404 33732 -12376
rect 33796 -12404 33852 -12376
rect 33916 -12404 33972 -12376
rect 34036 -12404 34092 -12376
rect 34156 -12404 34212 -12376
rect 34276 -12404 34332 -12376
rect 34396 -12404 34452 -12376
rect 34516 -12404 34572 -12376
rect 34636 -12404 34692 -12376
rect 34756 -12404 34812 -12376
rect 34876 -12404 34932 -12376
rect 34996 -12404 35052 -12376
rect 35116 -12404 35172 -12376
rect 35236 -12404 35292 -12376
rect 35356 -12404 35412 -12376
rect 35476 -12404 35532 -12376
rect 35596 -12404 35652 -12376
rect 35716 -12404 35772 -12376
rect 35836 -12404 35892 -12376
rect 35956 -12404 36012 -12376
rect 36076 -12404 36132 -12376
rect 36196 -12404 36252 -12376
rect 36316 -12404 36372 -12376
rect 36436 -12404 36492 -12376
rect 36556 -12404 36612 -12376
rect 36676 -12404 36732 -12376
rect 36796 -12404 36852 -12376
rect 36916 -12404 36972 -12376
rect 37036 -12404 37092 -12376
rect 37156 -12404 37212 -12376
rect 37276 -12404 37332 -12376
rect 37396 -12404 37452 -12376
rect 37516 -12404 37572 -12376
rect 37636 -12404 37692 -12376
rect 37756 -12404 37812 -12376
rect 37876 -12404 37932 -12376
rect 37996 -12404 38052 -12376
rect 38116 -12404 38172 -12376
rect 38236 -12404 38292 -12376
rect 38356 -12404 38412 -12376
rect 38476 -12404 38532 -12376
rect 38596 -12404 38652 -12376
rect 38716 -12404 38772 -12376
rect 38836 -12404 38892 -12376
rect 38956 -12404 39012 -12376
rect 39076 -12404 39132 -12376
rect 39196 -12404 39252 -12376
rect 39316 -12404 39372 -12376
rect 39436 -12404 39492 -12376
rect 39556 -12404 39612 -12376
rect 39676 -12404 39732 -12376
rect 39796 -12404 39852 -12376
rect 39916 -12404 39972 -12376
rect 40036 -12404 40092 -12376
rect 40156 -12404 40212 -12376
rect 40276 -12404 40332 -12376
rect 40396 -12404 40452 -12376
rect 40516 -12404 40572 -12376
rect 40636 -12404 40692 -12376
rect 40756 -12404 40812 -12376
rect 40876 -12404 40932 -12376
rect 40996 -12404 41052 -12376
rect 41116 -12404 41172 -12376
rect 41236 -12404 41292 -12376
rect 41356 -12404 41412 -12376
rect 41476 -12404 41532 -12376
rect 41596 -12404 41652 -12376
rect 41716 -12404 41772 -12376
rect 41836 -12404 41892 -12376
rect 41956 -12404 42012 -12376
rect 42076 -12404 42132 -12376
rect 42196 -12404 42252 -12376
rect 42316 -12404 42372 -12376
rect 42436 -12404 42492 -12376
rect 42556 -12404 42612 -12376
rect 42676 -12404 42732 -12376
rect 42796 -12404 42852 -12376
rect 42916 -12404 42972 -12376
rect 43036 -12404 43092 -12376
rect 43156 -12404 43212 -12376
rect 43276 -12404 43332 -12376
rect 43396 -12404 43452 -12376
rect 43516 -12404 43572 -12376
rect 43636 -12404 43692 -12376
rect 43756 -12404 43812 -12376
rect 43876 -12404 43932 -12376
rect 43996 -12404 44052 -12376
rect 44116 -12404 44172 -12376
rect 44236 -12404 44292 -12376
rect 44356 -12404 44412 -12376
rect 44476 -12404 44532 -12376
rect 44596 -12404 44652 -12376
rect 44716 -12404 44772 -12376
rect 44836 -12404 44892 -12376
rect 44956 -12404 45012 -12376
rect 45076 -12404 45132 -12376
rect 45196 -12404 45252 -12376
rect 45316 -12404 45372 -12376
rect 45436 -12404 45492 -12376
rect 45556 -12404 45612 -12376
rect 25848 -12548 25932 -12528
rect 25848 -12556 25868 -12548
rect 25876 -12556 25904 -12548
rect 25912 -12556 25932 -12548
rect 25968 -12548 26052 -12528
rect 25968 -12556 25988 -12548
rect 25996 -12556 26024 -12548
rect 26032 -12556 26052 -12548
rect 26088 -12548 26172 -12528
rect 26088 -12556 26108 -12548
rect 26116 -12556 26144 -12548
rect 26152 -12556 26172 -12548
rect 26208 -12548 26292 -12528
rect 26208 -12556 26228 -12548
rect 26236 -12556 26264 -12548
rect 26272 -12556 26292 -12548
rect 26328 -12548 26412 -12528
rect 26328 -12556 26348 -12548
rect 26356 -12556 26384 -12548
rect 26392 -12556 26412 -12548
rect 26448 -12548 26532 -12528
rect 26448 -12556 26468 -12548
rect 26476 -12556 26504 -12548
rect 26512 -12556 26532 -12548
rect 26568 -12548 26652 -12528
rect 26568 -12556 26588 -12548
rect 26596 -12556 26624 -12548
rect 26632 -12556 26652 -12548
rect 26688 -12548 26772 -12528
rect 26688 -12556 26708 -12548
rect 26716 -12556 26744 -12548
rect 26752 -12556 26772 -12548
rect 26808 -12548 26892 -12528
rect 26808 -12556 26828 -12548
rect 26836 -12556 26864 -12548
rect 26872 -12556 26892 -12548
rect 26928 -12548 27012 -12528
rect 26928 -12556 26948 -12548
rect 26956 -12556 26984 -12548
rect 26992 -12556 27012 -12548
rect 27048 -12548 27132 -12528
rect 27048 -12556 27068 -12548
rect 27076 -12556 27104 -12548
rect 27112 -12556 27132 -12548
rect 27168 -12548 27252 -12528
rect 27168 -12556 27188 -12548
rect 27196 -12556 27224 -12548
rect 27232 -12556 27252 -12548
rect 27288 -12548 27372 -12528
rect 27288 -12556 27308 -12548
rect 27316 -12556 27344 -12548
rect 27352 -12556 27372 -12548
rect 27408 -12548 27492 -12528
rect 27408 -12556 27428 -12548
rect 27436 -12556 27464 -12548
rect 27472 -12556 27492 -12548
rect 27528 -12548 27612 -12528
rect 27528 -12556 27548 -12548
rect 27556 -12556 27584 -12548
rect 27592 -12556 27612 -12548
rect 27648 -12548 27732 -12528
rect 27648 -12556 27668 -12548
rect 27676 -12556 27704 -12548
rect 27712 -12556 27732 -12548
rect 27768 -12548 27852 -12528
rect 27768 -12556 27788 -12548
rect 27796 -12556 27824 -12548
rect 27832 -12556 27852 -12548
rect 27888 -12548 27972 -12528
rect 27888 -12556 27908 -12548
rect 27916 -12556 27944 -12548
rect 27952 -12556 27972 -12548
rect 28008 -12548 28092 -12528
rect 28008 -12556 28028 -12548
rect 28036 -12556 28064 -12548
rect 28072 -12556 28092 -12548
rect 28128 -12548 28212 -12528
rect 28128 -12556 28148 -12548
rect 28156 -12556 28184 -12548
rect 28192 -12556 28212 -12548
rect 28248 -12548 28332 -12528
rect 28248 -12556 28268 -12548
rect 28276 -12556 28304 -12548
rect 28312 -12556 28332 -12548
rect 28368 -12548 28452 -12528
rect 28368 -12556 28388 -12548
rect 28396 -12556 28424 -12548
rect 28432 -12556 28452 -12548
rect 28488 -12548 28572 -12528
rect 28488 -12556 28508 -12548
rect 28516 -12556 28544 -12548
rect 28552 -12556 28572 -12548
rect 28608 -12548 28692 -12528
rect 28608 -12556 28628 -12548
rect 28636 -12556 28664 -12548
rect 28672 -12556 28692 -12548
rect 28728 -12548 28812 -12528
rect 28728 -12556 28748 -12548
rect 28756 -12556 28784 -12548
rect 28792 -12556 28812 -12548
rect 28848 -12548 28932 -12528
rect 28848 -12556 28868 -12548
rect 28876 -12556 28904 -12548
rect 28912 -12556 28932 -12548
rect 28968 -12548 29052 -12528
rect 28968 -12556 28988 -12548
rect 28996 -12556 29024 -12548
rect 29032 -12556 29052 -12548
rect 29088 -12548 29172 -12528
rect 29088 -12556 29108 -12548
rect 29116 -12556 29144 -12548
rect 29152 -12556 29172 -12548
rect 29208 -12548 29292 -12528
rect 29208 -12556 29228 -12548
rect 29236 -12556 29264 -12548
rect 29272 -12556 29292 -12548
rect 29328 -12548 29412 -12528
rect 29328 -12556 29348 -12548
rect 29356 -12556 29384 -12548
rect 29392 -12556 29412 -12548
rect 29448 -12548 29532 -12528
rect 29448 -12556 29468 -12548
rect 29476 -12556 29504 -12548
rect 29512 -12556 29532 -12548
rect 29568 -12548 29652 -12528
rect 29568 -12556 29588 -12548
rect 29596 -12556 29624 -12548
rect 29632 -12556 29652 -12548
rect 29688 -12548 29772 -12528
rect 29688 -12556 29708 -12548
rect 29716 -12556 29744 -12548
rect 29752 -12556 29772 -12548
rect 29808 -12548 29892 -12528
rect 29808 -12556 29828 -12548
rect 29836 -12556 29864 -12548
rect 29872 -12556 29892 -12548
rect 29928 -12548 30012 -12528
rect 29928 -12556 29948 -12548
rect 29956 -12556 29984 -12548
rect 29992 -12556 30012 -12548
rect 30048 -12548 30132 -12528
rect 30048 -12556 30068 -12548
rect 30076 -12556 30104 -12548
rect 30112 -12556 30132 -12548
rect 30168 -12548 30252 -12528
rect 30168 -12556 30188 -12548
rect 30196 -12556 30224 -12548
rect 30232 -12556 30252 -12548
rect 30288 -12548 30372 -12528
rect 30288 -12556 30308 -12548
rect 30316 -12556 30344 -12548
rect 30352 -12556 30372 -12548
rect 30408 -12548 30492 -12528
rect 30408 -12556 30428 -12548
rect 30436 -12556 30464 -12548
rect 30472 -12556 30492 -12548
rect 30528 -12548 30612 -12528
rect 30528 -12556 30548 -12548
rect 30556 -12556 30584 -12548
rect 30592 -12556 30612 -12548
rect 30648 -12548 30732 -12528
rect 30648 -12556 30668 -12548
rect 30676 -12556 30704 -12548
rect 30712 -12556 30732 -12548
rect 30768 -12548 30852 -12528
rect 30768 -12556 30788 -12548
rect 30796 -12556 30824 -12548
rect 30832 -12556 30852 -12548
rect 30888 -12548 30972 -12528
rect 30888 -12556 30908 -12548
rect 30916 -12556 30944 -12548
rect 30952 -12556 30972 -12548
rect 31008 -12548 31092 -12528
rect 31008 -12556 31028 -12548
rect 31036 -12556 31064 -12548
rect 31072 -12556 31092 -12548
rect 31128 -12548 31212 -12528
rect 31128 -12556 31148 -12548
rect 31156 -12556 31184 -12548
rect 31192 -12556 31212 -12548
rect 31248 -12548 31332 -12528
rect 31248 -12556 31268 -12548
rect 31276 -12556 31304 -12548
rect 31312 -12556 31332 -12548
rect 31368 -12548 31452 -12528
rect 31368 -12556 31388 -12548
rect 31396 -12556 31424 -12548
rect 31432 -12556 31452 -12548
rect 31488 -12548 31572 -12528
rect 31488 -12556 31508 -12548
rect 31516 -12556 31544 -12548
rect 31552 -12556 31572 -12548
rect 31608 -12548 31692 -12528
rect 31608 -12556 31628 -12548
rect 31636 -12556 31664 -12548
rect 31672 -12556 31692 -12548
rect 31728 -12548 31812 -12528
rect 31728 -12556 31748 -12548
rect 31756 -12556 31784 -12548
rect 31792 -12556 31812 -12548
rect 31848 -12548 31932 -12528
rect 31848 -12556 31868 -12548
rect 31876 -12556 31904 -12548
rect 31912 -12556 31932 -12548
rect 31968 -12548 32052 -12528
rect 31968 -12556 31988 -12548
rect 31996 -12556 32024 -12548
rect 32032 -12556 32052 -12548
rect 32088 -12548 32172 -12528
rect 32088 -12556 32108 -12548
rect 32116 -12556 32144 -12548
rect 32152 -12556 32172 -12548
rect 32208 -12548 32292 -12528
rect 32208 -12556 32228 -12548
rect 32236 -12556 32264 -12548
rect 32272 -12556 32292 -12548
rect 32328 -12548 32412 -12528
rect 32328 -12556 32348 -12548
rect 32356 -12556 32384 -12548
rect 32392 -12556 32412 -12548
rect 32448 -12548 32532 -12528
rect 32448 -12556 32468 -12548
rect 32476 -12556 32504 -12548
rect 32512 -12556 32532 -12548
rect 32568 -12548 32652 -12528
rect 32568 -12556 32588 -12548
rect 32596 -12556 32624 -12548
rect 32632 -12556 32652 -12548
rect 32688 -12548 32772 -12528
rect 32688 -12556 32708 -12548
rect 32716 -12556 32744 -12548
rect 32752 -12556 32772 -12548
rect 32808 -12548 32892 -12528
rect 32808 -12556 32828 -12548
rect 32836 -12556 32864 -12548
rect 32872 -12556 32892 -12548
rect 32928 -12548 33012 -12528
rect 32928 -12556 32948 -12548
rect 32956 -12556 32984 -12548
rect 32992 -12556 33012 -12548
rect 33048 -12548 33132 -12528
rect 33048 -12556 33068 -12548
rect 33076 -12556 33104 -12548
rect 33112 -12556 33132 -12548
rect 33168 -12548 33252 -12528
rect 33168 -12556 33188 -12548
rect 33196 -12556 33224 -12548
rect 33232 -12556 33252 -12548
rect 33288 -12548 33372 -12528
rect 33288 -12556 33308 -12548
rect 33316 -12556 33344 -12548
rect 33352 -12556 33372 -12548
rect 33408 -12548 33492 -12528
rect 33408 -12556 33428 -12548
rect 33436 -12556 33464 -12548
rect 33472 -12556 33492 -12548
rect 33528 -12548 33612 -12528
rect 33528 -12556 33548 -12548
rect 33556 -12556 33584 -12548
rect 33592 -12556 33612 -12548
rect 33648 -12548 33732 -12528
rect 33648 -12556 33668 -12548
rect 33676 -12556 33704 -12548
rect 33712 -12556 33732 -12548
rect 33768 -12548 33852 -12528
rect 33768 -12556 33788 -12548
rect 33796 -12556 33824 -12548
rect 33832 -12556 33852 -12548
rect 33888 -12548 33972 -12528
rect 33888 -12556 33908 -12548
rect 33916 -12556 33944 -12548
rect 33952 -12556 33972 -12548
rect 34008 -12548 34092 -12528
rect 34008 -12556 34028 -12548
rect 34036 -12556 34064 -12548
rect 34072 -12556 34092 -12548
rect 34128 -12548 34212 -12528
rect 34128 -12556 34148 -12548
rect 34156 -12556 34184 -12548
rect 34192 -12556 34212 -12548
rect 34248 -12548 34332 -12528
rect 34248 -12556 34268 -12548
rect 34276 -12556 34304 -12548
rect 34312 -12556 34332 -12548
rect 34368 -12548 34452 -12528
rect 34368 -12556 34388 -12548
rect 34396 -12556 34424 -12548
rect 34432 -12556 34452 -12548
rect 34488 -12548 34572 -12528
rect 34488 -12556 34508 -12548
rect 34516 -12556 34544 -12548
rect 34552 -12556 34572 -12548
rect 34608 -12548 34692 -12528
rect 34608 -12556 34628 -12548
rect 34636 -12556 34664 -12548
rect 34672 -12556 34692 -12548
rect 34728 -12548 34812 -12528
rect 34728 -12556 34748 -12548
rect 34756 -12556 34784 -12548
rect 34792 -12556 34812 -12548
rect 34848 -12548 34932 -12528
rect 34848 -12556 34868 -12548
rect 34876 -12556 34904 -12548
rect 34912 -12556 34932 -12548
rect 34968 -12548 35052 -12528
rect 34968 -12556 34988 -12548
rect 34996 -12556 35024 -12548
rect 35032 -12556 35052 -12548
rect 35088 -12548 35172 -12528
rect 35088 -12556 35108 -12548
rect 35116 -12556 35144 -12548
rect 35152 -12556 35172 -12548
rect 35208 -12548 35292 -12528
rect 35208 -12556 35228 -12548
rect 35236 -12556 35264 -12548
rect 35272 -12556 35292 -12548
rect 35328 -12548 35412 -12528
rect 35328 -12556 35348 -12548
rect 35356 -12556 35384 -12548
rect 35392 -12556 35412 -12548
rect 35448 -12548 35532 -12528
rect 35448 -12556 35468 -12548
rect 35476 -12556 35504 -12548
rect 35512 -12556 35532 -12548
rect 35568 -12548 35652 -12528
rect 35568 -12556 35588 -12548
rect 35596 -12556 35624 -12548
rect 35632 -12556 35652 -12548
rect 35688 -12548 35772 -12528
rect 35688 -12556 35708 -12548
rect 35716 -12556 35744 -12548
rect 35752 -12556 35772 -12548
rect 35808 -12548 35892 -12528
rect 35808 -12556 35828 -12548
rect 35836 -12556 35864 -12548
rect 35872 -12556 35892 -12548
rect 35928 -12548 36012 -12528
rect 35928 -12556 35948 -12548
rect 35956 -12556 35984 -12548
rect 35992 -12556 36012 -12548
rect 36048 -12548 36132 -12528
rect 36048 -12556 36068 -12548
rect 36076 -12556 36104 -12548
rect 36112 -12556 36132 -12548
rect 36168 -12548 36252 -12528
rect 36168 -12556 36188 -12548
rect 36196 -12556 36224 -12548
rect 36232 -12556 36252 -12548
rect 36288 -12548 36372 -12528
rect 36288 -12556 36308 -12548
rect 36316 -12556 36344 -12548
rect 36352 -12556 36372 -12548
rect 36408 -12548 36492 -12528
rect 36408 -12556 36428 -12548
rect 36436 -12556 36464 -12548
rect 36472 -12556 36492 -12548
rect 36528 -12548 36612 -12528
rect 36528 -12556 36548 -12548
rect 36556 -12556 36584 -12548
rect 36592 -12556 36612 -12548
rect 36648 -12548 36732 -12528
rect 36648 -12556 36668 -12548
rect 36676 -12556 36704 -12548
rect 36712 -12556 36732 -12548
rect 36768 -12548 36852 -12528
rect 36768 -12556 36788 -12548
rect 36796 -12556 36824 -12548
rect 36832 -12556 36852 -12548
rect 36888 -12548 36972 -12528
rect 36888 -12556 36908 -12548
rect 36916 -12556 36944 -12548
rect 36952 -12556 36972 -12548
rect 37008 -12548 37092 -12528
rect 37008 -12556 37028 -12548
rect 37036 -12556 37064 -12548
rect 37072 -12556 37092 -12548
rect 37128 -12548 37212 -12528
rect 37128 -12556 37148 -12548
rect 37156 -12556 37184 -12548
rect 37192 -12556 37212 -12548
rect 37248 -12548 37332 -12528
rect 37248 -12556 37268 -12548
rect 37276 -12556 37304 -12548
rect 37312 -12556 37332 -12548
rect 37368 -12548 37452 -12528
rect 37368 -12556 37388 -12548
rect 37396 -12556 37424 -12548
rect 37432 -12556 37452 -12548
rect 37488 -12548 37572 -12528
rect 37488 -12556 37508 -12548
rect 37516 -12556 37544 -12548
rect 37552 -12556 37572 -12548
rect 37608 -12548 37692 -12528
rect 37608 -12556 37628 -12548
rect 37636 -12556 37664 -12548
rect 37672 -12556 37692 -12548
rect 37728 -12548 37812 -12528
rect 37728 -12556 37748 -12548
rect 37756 -12556 37784 -12548
rect 37792 -12556 37812 -12548
rect 37848 -12548 37932 -12528
rect 37848 -12556 37868 -12548
rect 37876 -12556 37904 -12548
rect 37912 -12556 37932 -12548
rect 37968 -12548 38052 -12528
rect 37968 -12556 37988 -12548
rect 37996 -12556 38024 -12548
rect 38032 -12556 38052 -12548
rect 38088 -12548 38172 -12528
rect 38088 -12556 38108 -12548
rect 38116 -12556 38144 -12548
rect 38152 -12556 38172 -12548
rect 38208 -12548 38292 -12528
rect 38208 -12556 38228 -12548
rect 38236 -12556 38264 -12548
rect 38272 -12556 38292 -12548
rect 38328 -12548 38412 -12528
rect 38328 -12556 38348 -12548
rect 38356 -12556 38384 -12548
rect 38392 -12556 38412 -12548
rect 38448 -12548 38532 -12528
rect 38448 -12556 38468 -12548
rect 38476 -12556 38504 -12548
rect 38512 -12556 38532 -12548
rect 38568 -12548 38652 -12528
rect 38568 -12556 38588 -12548
rect 38596 -12556 38624 -12548
rect 38632 -12556 38652 -12548
rect 38688 -12548 38772 -12528
rect 38688 -12556 38708 -12548
rect 38716 -12556 38744 -12548
rect 38752 -12556 38772 -12548
rect 38808 -12548 38892 -12528
rect 38808 -12556 38828 -12548
rect 38836 -12556 38864 -12548
rect 38872 -12556 38892 -12548
rect 38928 -12548 39012 -12528
rect 38928 -12556 38948 -12548
rect 38956 -12556 38984 -12548
rect 38992 -12556 39012 -12548
rect 39048 -12548 39132 -12528
rect 39048 -12556 39068 -12548
rect 39076 -12556 39104 -12548
rect 39112 -12556 39132 -12548
rect 39168 -12548 39252 -12528
rect 39168 -12556 39188 -12548
rect 39196 -12556 39224 -12548
rect 39232 -12556 39252 -12548
rect 39288 -12548 39372 -12528
rect 39288 -12556 39308 -12548
rect 39316 -12556 39344 -12548
rect 39352 -12556 39372 -12548
rect 39408 -12548 39492 -12528
rect 39408 -12556 39428 -12548
rect 39436 -12556 39464 -12548
rect 39472 -12556 39492 -12548
rect 39528 -12548 39612 -12528
rect 39528 -12556 39548 -12548
rect 39556 -12556 39584 -12548
rect 39592 -12556 39612 -12548
rect 39648 -12548 39732 -12528
rect 39648 -12556 39668 -12548
rect 39676 -12556 39704 -12548
rect 39712 -12556 39732 -12548
rect 39768 -12548 39852 -12528
rect 39768 -12556 39788 -12548
rect 39796 -12556 39824 -12548
rect 39832 -12556 39852 -12548
rect 39888 -12548 39972 -12528
rect 39888 -12556 39908 -12548
rect 39916 -12556 39944 -12548
rect 39952 -12556 39972 -12548
rect 40008 -12548 40092 -12528
rect 40008 -12556 40028 -12548
rect 40036 -12556 40064 -12548
rect 40072 -12556 40092 -12548
rect 40128 -12548 40212 -12528
rect 40128 -12556 40148 -12548
rect 40156 -12556 40184 -12548
rect 40192 -12556 40212 -12548
rect 40248 -12548 40332 -12528
rect 40248 -12556 40268 -12548
rect 40276 -12556 40304 -12548
rect 40312 -12556 40332 -12548
rect 40368 -12548 40452 -12528
rect 40368 -12556 40388 -12548
rect 40396 -12556 40424 -12548
rect 40432 -12556 40452 -12548
rect 40488 -12548 40572 -12528
rect 40488 -12556 40508 -12548
rect 40516 -12556 40544 -12548
rect 40552 -12556 40572 -12548
rect 40608 -12548 40692 -12528
rect 40608 -12556 40628 -12548
rect 40636 -12556 40664 -12548
rect 40672 -12556 40692 -12548
rect 40728 -12548 40812 -12528
rect 40728 -12556 40748 -12548
rect 40756 -12556 40784 -12548
rect 40792 -12556 40812 -12548
rect 40848 -12548 40932 -12528
rect 40848 -12556 40868 -12548
rect 40876 -12556 40904 -12548
rect 40912 -12556 40932 -12548
rect 40968 -12548 41052 -12528
rect 40968 -12556 40988 -12548
rect 40996 -12556 41024 -12548
rect 41032 -12556 41052 -12548
rect 41088 -12548 41172 -12528
rect 41088 -12556 41108 -12548
rect 41116 -12556 41144 -12548
rect 41152 -12556 41172 -12548
rect 41208 -12548 41292 -12528
rect 41208 -12556 41228 -12548
rect 41236 -12556 41264 -12548
rect 41272 -12556 41292 -12548
rect 41328 -12548 41412 -12528
rect 41328 -12556 41348 -12548
rect 41356 -12556 41384 -12548
rect 41392 -12556 41412 -12548
rect 41448 -12548 41532 -12528
rect 41448 -12556 41468 -12548
rect 41476 -12556 41504 -12548
rect 41512 -12556 41532 -12548
rect 41568 -12548 41652 -12528
rect 41568 -12556 41588 -12548
rect 41596 -12556 41624 -12548
rect 41632 -12556 41652 -12548
rect 41688 -12548 41772 -12528
rect 41688 -12556 41708 -12548
rect 41716 -12556 41744 -12548
rect 41752 -12556 41772 -12548
rect 41808 -12548 41892 -12528
rect 41808 -12556 41828 -12548
rect 41836 -12556 41864 -12548
rect 41872 -12556 41892 -12548
rect 41928 -12548 42012 -12528
rect 41928 -12556 41948 -12548
rect 41956 -12556 41984 -12548
rect 41992 -12556 42012 -12548
rect 42048 -12548 42132 -12528
rect 42048 -12556 42068 -12548
rect 42076 -12556 42104 -12548
rect 42112 -12556 42132 -12548
rect 42168 -12548 42252 -12528
rect 42168 -12556 42188 -12548
rect 42196 -12556 42224 -12548
rect 42232 -12556 42252 -12548
rect 42288 -12548 42372 -12528
rect 42288 -12556 42308 -12548
rect 42316 -12556 42344 -12548
rect 42352 -12556 42372 -12548
rect 42408 -12548 42492 -12528
rect 42408 -12556 42428 -12548
rect 42436 -12556 42464 -12548
rect 42472 -12556 42492 -12548
rect 42528 -12548 42612 -12528
rect 42528 -12556 42548 -12548
rect 42556 -12556 42584 -12548
rect 42592 -12556 42612 -12548
rect 42648 -12548 42732 -12528
rect 42648 -12556 42668 -12548
rect 42676 -12556 42704 -12548
rect 42712 -12556 42732 -12548
rect 42768 -12548 42852 -12528
rect 42768 -12556 42788 -12548
rect 42796 -12556 42824 -12548
rect 42832 -12556 42852 -12548
rect 42888 -12548 42972 -12528
rect 42888 -12556 42908 -12548
rect 42916 -12556 42944 -12548
rect 42952 -12556 42972 -12548
rect 43008 -12548 43092 -12528
rect 43008 -12556 43028 -12548
rect 43036 -12556 43064 -12548
rect 43072 -12556 43092 -12548
rect 43128 -12548 43212 -12528
rect 43128 -12556 43148 -12548
rect 43156 -12556 43184 -12548
rect 43192 -12556 43212 -12548
rect 43248 -12548 43332 -12528
rect 43248 -12556 43268 -12548
rect 43276 -12556 43304 -12548
rect 43312 -12556 43332 -12548
rect 43368 -12548 43452 -12528
rect 43368 -12556 43388 -12548
rect 43396 -12556 43424 -12548
rect 43432 -12556 43452 -12548
rect 43488 -12548 43572 -12528
rect 43488 -12556 43508 -12548
rect 43516 -12556 43544 -12548
rect 43552 -12556 43572 -12548
rect 43608 -12548 43692 -12528
rect 43608 -12556 43628 -12548
rect 43636 -12556 43664 -12548
rect 43672 -12556 43692 -12548
rect 43728 -12548 43812 -12528
rect 43728 -12556 43748 -12548
rect 43756 -12556 43784 -12548
rect 43792 -12556 43812 -12548
rect 43848 -12548 43932 -12528
rect 43848 -12556 43868 -12548
rect 43876 -12556 43904 -12548
rect 43912 -12556 43932 -12548
rect 43968 -12548 44052 -12528
rect 43968 -12556 43988 -12548
rect 43996 -12556 44024 -12548
rect 44032 -12556 44052 -12548
rect 44088 -12548 44172 -12528
rect 44088 -12556 44108 -12548
rect 44116 -12556 44144 -12548
rect 44152 -12556 44172 -12548
rect 44208 -12548 44292 -12528
rect 44208 -12556 44228 -12548
rect 44236 -12556 44264 -12548
rect 44272 -12556 44292 -12548
rect 44328 -12548 44412 -12528
rect 44328 -12556 44348 -12548
rect 44356 -12556 44384 -12548
rect 44392 -12556 44412 -12548
rect 44448 -12548 44532 -12528
rect 44448 -12556 44468 -12548
rect 44476 -12556 44504 -12548
rect 44512 -12556 44532 -12548
rect 44568 -12548 44652 -12528
rect 44568 -12556 44588 -12548
rect 44596 -12556 44624 -12548
rect 44632 -12556 44652 -12548
rect 44688 -12548 44772 -12528
rect 44688 -12556 44708 -12548
rect 44716 -12556 44744 -12548
rect 44752 -12556 44772 -12548
rect 44808 -12548 44892 -12528
rect 44808 -12556 44828 -12548
rect 44836 -12556 44864 -12548
rect 44872 -12556 44892 -12548
rect 44928 -12548 45012 -12528
rect 44928 -12556 44948 -12548
rect 44956 -12556 44984 -12548
rect 44992 -12556 45012 -12548
rect 45048 -12548 45132 -12528
rect 45048 -12556 45068 -12548
rect 45076 -12556 45104 -12548
rect 45112 -12556 45132 -12548
rect 45168 -12548 45252 -12528
rect 45168 -12556 45188 -12548
rect 45196 -12556 45224 -12548
rect 45232 -12556 45252 -12548
rect 45288 -12548 45372 -12528
rect 45288 -12556 45308 -12548
rect 45316 -12556 45344 -12548
rect 45352 -12556 45372 -12548
rect 45408 -12548 45492 -12528
rect 45408 -12556 45428 -12548
rect 45436 -12556 45464 -12548
rect 45472 -12556 45492 -12548
rect 45528 -12548 45612 -12528
rect 45528 -12556 45548 -12548
rect 45556 -12556 45584 -12548
rect 45592 -12556 45612 -12548
rect 25876 -12584 25932 -12556
rect 25996 -12584 26052 -12556
rect 26116 -12584 26172 -12556
rect 26236 -12584 26292 -12556
rect 26356 -12584 26412 -12556
rect 26476 -12584 26532 -12556
rect 26596 -12584 26652 -12556
rect 26716 -12584 26772 -12556
rect 26836 -12584 26892 -12556
rect 26956 -12584 27012 -12556
rect 27076 -12584 27132 -12556
rect 27196 -12584 27252 -12556
rect 27316 -12584 27372 -12556
rect 27436 -12584 27492 -12556
rect 27556 -12584 27612 -12556
rect 27676 -12584 27732 -12556
rect 27796 -12584 27852 -12556
rect 27916 -12584 27972 -12556
rect 28036 -12584 28092 -12556
rect 28156 -12584 28212 -12556
rect 28276 -12584 28332 -12556
rect 28396 -12584 28452 -12556
rect 28516 -12584 28572 -12556
rect 28636 -12584 28692 -12556
rect 28756 -12584 28812 -12556
rect 28876 -12584 28932 -12556
rect 28996 -12584 29052 -12556
rect 29116 -12584 29172 -12556
rect 29236 -12584 29292 -12556
rect 29356 -12584 29412 -12556
rect 29476 -12584 29532 -12556
rect 29596 -12584 29652 -12556
rect 29716 -12584 29772 -12556
rect 29836 -12584 29892 -12556
rect 29956 -12584 30012 -12556
rect 30076 -12584 30132 -12556
rect 30196 -12584 30252 -12556
rect 30316 -12584 30372 -12556
rect 30436 -12584 30492 -12556
rect 30556 -12584 30612 -12556
rect 30676 -12584 30732 -12556
rect 30796 -12584 30852 -12556
rect 30916 -12584 30972 -12556
rect 31036 -12584 31092 -12556
rect 31156 -12584 31212 -12556
rect 31276 -12584 31332 -12556
rect 31396 -12584 31452 -12556
rect 31516 -12584 31572 -12556
rect 31636 -12584 31692 -12556
rect 31756 -12584 31812 -12556
rect 31876 -12584 31932 -12556
rect 31996 -12584 32052 -12556
rect 32116 -12584 32172 -12556
rect 32236 -12584 32292 -12556
rect 32356 -12584 32412 -12556
rect 32476 -12584 32532 -12556
rect 32596 -12584 32652 -12556
rect 32716 -12584 32772 -12556
rect 32836 -12584 32892 -12556
rect 32956 -12584 33012 -12556
rect 33076 -12584 33132 -12556
rect 33196 -12584 33252 -12556
rect 33316 -12584 33372 -12556
rect 33436 -12584 33492 -12556
rect 33556 -12584 33612 -12556
rect 33676 -12584 33732 -12556
rect 33796 -12584 33852 -12556
rect 33916 -12584 33972 -12556
rect 34036 -12584 34092 -12556
rect 34156 -12584 34212 -12556
rect 34276 -12584 34332 -12556
rect 34396 -12584 34452 -12556
rect 34516 -12584 34572 -12556
rect 34636 -12584 34692 -12556
rect 34756 -12584 34812 -12556
rect 34876 -12584 34932 -12556
rect 34996 -12584 35052 -12556
rect 35116 -12584 35172 -12556
rect 35236 -12584 35292 -12556
rect 35356 -12584 35412 -12556
rect 35476 -12584 35532 -12556
rect 35596 -12584 35652 -12556
rect 35716 -12584 35772 -12556
rect 35836 -12584 35892 -12556
rect 35956 -12584 36012 -12556
rect 36076 -12584 36132 -12556
rect 36196 -12584 36252 -12556
rect 36316 -12584 36372 -12556
rect 36436 -12584 36492 -12556
rect 36556 -12584 36612 -12556
rect 36676 -12584 36732 -12556
rect 36796 -12584 36852 -12556
rect 36916 -12584 36972 -12556
rect 37036 -12584 37092 -12556
rect 37156 -12584 37212 -12556
rect 37276 -12584 37332 -12556
rect 37396 -12584 37452 -12556
rect 37516 -12584 37572 -12556
rect 37636 -12584 37692 -12556
rect 37756 -12584 37812 -12556
rect 37876 -12584 37932 -12556
rect 37996 -12584 38052 -12556
rect 38116 -12584 38172 -12556
rect 38236 -12584 38292 -12556
rect 38356 -12584 38412 -12556
rect 38476 -12584 38532 -12556
rect 38596 -12584 38652 -12556
rect 38716 -12584 38772 -12556
rect 38836 -12584 38892 -12556
rect 38956 -12584 39012 -12556
rect 39076 -12584 39132 -12556
rect 39196 -12584 39252 -12556
rect 39316 -12584 39372 -12556
rect 39436 -12584 39492 -12556
rect 39556 -12584 39612 -12556
rect 39676 -12584 39732 -12556
rect 39796 -12584 39852 -12556
rect 39916 -12584 39972 -12556
rect 40036 -12584 40092 -12556
rect 40156 -12584 40212 -12556
rect 40276 -12584 40332 -12556
rect 40396 -12584 40452 -12556
rect 40516 -12584 40572 -12556
rect 40636 -12584 40692 -12556
rect 40756 -12584 40812 -12556
rect 40876 -12584 40932 -12556
rect 40996 -12584 41052 -12556
rect 41116 -12584 41172 -12556
rect 41236 -12584 41292 -12556
rect 41356 -12584 41412 -12556
rect 41476 -12584 41532 -12556
rect 41596 -12584 41652 -12556
rect 41716 -12584 41772 -12556
rect 41836 -12584 41892 -12556
rect 41956 -12584 42012 -12556
rect 42076 -12584 42132 -12556
rect 42196 -12584 42252 -12556
rect 42316 -12584 42372 -12556
rect 42436 -12584 42492 -12556
rect 42556 -12584 42612 -12556
rect 42676 -12584 42732 -12556
rect 42796 -12584 42852 -12556
rect 42916 -12584 42972 -12556
rect 43036 -12584 43092 -12556
rect 43156 -12584 43212 -12556
rect 43276 -12584 43332 -12556
rect 43396 -12584 43452 -12556
rect 43516 -12584 43572 -12556
rect 43636 -12584 43692 -12556
rect 43756 -12584 43812 -12556
rect 43876 -12584 43932 -12556
rect 43996 -12584 44052 -12556
rect 44116 -12584 44172 -12556
rect 44236 -12584 44292 -12556
rect 44356 -12584 44412 -12556
rect 44476 -12584 44532 -12556
rect 44596 -12584 44652 -12556
rect 44716 -12584 44772 -12556
rect 44836 -12584 44892 -12556
rect 44956 -12584 45012 -12556
rect 45076 -12584 45132 -12556
rect 45196 -12584 45252 -12556
rect 45316 -12584 45372 -12556
rect 45436 -12584 45492 -12556
rect 45556 -12584 45612 -12556
use barth_a  barth_a_0
timestamp 1663412335
transform 1 0 6960 0 1 -3060
box -5220 -840 2940 2880
use barthmanf_a  barthmanf_a_0
timestamp 1665148219
transform 1 0 16980 0 1 -10440
box -4680 -900 7080 3060
use barthnauta_a  barthnauta_a_0
timestamp 1663414815
transform 1 0 17520 0 1 -3060
box -5220 -840 5340 2880
use manf_a  manf_a_0
timestamp 1665149341
transform 1 0 6420 0 1 -10440
box -4680 -900 4680 3060
use manfvieru_a  manfvieru_a_0
timestamp 1665299032
transform 1 0 30840 0 1 -10740
box -5580 -1980 16140 4500
use nauta  nauta_0
timestamp 1665184495
transform 1 0 7020 0 1 4380
box -5220 -840 540 2640
use nautanauta_a  nautanauta_a_0
timestamp 1665298770
transform 1 0 30900 0 1 4380
box -5580 -1980 14940 4080
use nautavieru_a  nautavieru_a_0
timestamp 1665298688
transform 1 0 30840 0 1 -3060
box -5580 -1980 14940 4260
<< end >>
