magic
tech gf180mcuC
magscale 1 5
timestamp 1665184495
<< metal2 >>
rect -3900 1434 -3840 1440
rect -3900 1146 -3884 1434
rect -3856 1146 -3840 1434
rect -3900 1140 -3840 1146
rect -300 1434 -240 1440
rect -300 1146 -284 1434
rect -256 1146 -240 1434
rect -300 1140 -240 1146
rect 300 1434 360 1440
rect 300 1146 316 1434
rect 344 1146 360 1434
rect 300 1140 360 1146
rect 3900 1434 3960 1440
rect 3900 1146 3916 1434
rect 3944 1146 3960 1434
rect 3900 1140 3960 1146
rect -2700 704 -2640 720
rect -2700 676 -2684 704
rect -2656 676 -2640 704
rect -2700 660 -2640 676
rect -2100 704 -2040 720
rect -2100 676 -2084 704
rect -2056 676 -2040 704
rect -2100 660 -2040 676
rect 2100 704 2160 720
rect 2100 676 2116 704
rect 2144 676 2160 704
rect 2100 660 2160 676
rect 2700 704 2760 720
rect 2700 676 2716 704
rect 2744 676 2760 704
rect 2700 660 2760 676
rect -1500 464 -1440 480
rect -1500 436 -1484 464
rect -1456 436 -1440 464
rect -1500 420 -1440 436
rect 1500 464 1560 480
rect 1500 436 1516 464
rect 1544 436 1560 464
rect 1500 420 1560 436
rect -3300 -6 -3240 0
rect -3300 -294 -3284 -6
rect -3256 -294 -3240 -6
rect -3300 -300 -3240 -294
rect -900 -6 -840 0
rect -900 -294 -884 -6
rect -856 -294 -840 -6
rect -900 -300 -840 -294
rect 900 -6 960 0
rect 900 -294 916 -6
rect 944 -294 960 -6
rect 900 -300 960 -294
rect 3300 -6 3360 0
rect 3300 -294 3316 -6
rect 3344 -294 3360 -6
rect 3300 -300 3360 -294
<< via2 >>
rect -3884 1146 -3856 1434
rect -284 1146 -256 1434
rect 316 1146 344 1434
rect 3916 1146 3944 1434
rect -2684 676 -2656 704
rect -2084 676 -2056 704
rect 2116 676 2144 704
rect 2716 676 2744 704
rect -1484 436 -1456 464
rect 1516 436 1544 464
rect -3284 -294 -3256 -6
rect -884 -294 -856 -6
rect 916 -294 944 -6
rect 3316 -294 3344 -6
<< metal3 >>
rect -4680 2640 -4620 2940
rect -4680 2400 -4620 2460
rect -4680 2280 -4620 2340
rect -4680 1620 -4620 1680
rect -4680 1140 -4620 1440
rect -3900 1434 -3840 1440
rect -3900 1146 -3884 1434
rect -3856 1146 -3840 1434
rect -3900 1140 -3840 1146
rect -1980 1434 -1920 1440
rect -1980 1146 -1964 1434
rect -1936 1146 -1920 1434
rect -1980 1140 -1920 1146
rect -300 1434 -240 1440
rect -300 1146 -284 1434
rect -256 1146 -240 1434
rect -300 1140 -240 1146
rect 300 1434 360 1440
rect 300 1146 316 1434
rect 344 1146 360 1434
rect 300 1140 360 1146
rect 1980 1434 2040 1440
rect 1980 1146 1996 1434
rect 2024 1146 2040 1434
rect 1980 1140 2040 1146
rect 3900 1434 3960 1440
rect 3900 1146 3916 1434
rect 3944 1146 3960 1434
rect 3900 1140 3960 1146
rect -4680 900 -4620 960
rect -4020 944 -3960 960
rect -4020 916 -4004 944
rect -3976 916 -3960 944
rect -4020 900 -3960 916
rect -180 944 -120 960
rect -180 916 -164 944
rect -136 916 -120 944
rect -180 900 -120 916
rect 180 944 240 960
rect 180 916 196 944
rect 224 916 240 944
rect 180 900 240 916
rect 4020 944 4080 960
rect 4020 916 4036 944
rect 4064 916 4080 944
rect 4020 900 4080 916
rect -4680 660 -4620 720
rect -2700 704 -2640 720
rect -2700 676 -2684 704
rect -2656 676 -2640 704
rect -2700 660 -2640 676
rect -2580 704 -2520 720
rect -2580 676 -2564 704
rect -2536 676 -2520 704
rect -2580 660 -2520 676
rect -2220 704 -2160 720
rect -2220 676 -2204 704
rect -2176 676 -2160 704
rect -2220 660 -2160 676
rect -2100 704 -2040 720
rect -2100 676 -2084 704
rect -2056 676 -2040 704
rect -2100 660 -2040 676
rect -1620 704 -1560 720
rect -1620 676 -1604 704
rect -1576 676 -1560 704
rect -1620 660 -1560 676
rect 1620 704 1680 720
rect 1620 676 1636 704
rect 1664 676 1680 704
rect 1620 660 1680 676
rect 2100 704 2160 720
rect 2100 676 2116 704
rect 2144 676 2160 704
rect 2100 660 2160 676
rect 2220 704 2280 720
rect 2220 676 2236 704
rect 2264 676 2280 704
rect 2220 660 2280 676
rect 2580 704 2640 720
rect 2580 676 2596 704
rect 2624 676 2640 704
rect 2580 660 2640 676
rect 2700 704 2760 720
rect 2700 676 2716 704
rect 2744 676 2760 704
rect 2700 660 2760 676
rect -4680 420 -4620 480
rect -3780 464 -3720 480
rect -3780 436 -3764 464
rect -3736 436 -3720 464
rect -3780 420 -3720 436
rect -3420 464 -3360 480
rect -3420 436 -3404 464
rect -3376 436 -3360 464
rect -3420 420 -3360 436
rect -1500 464 -1440 480
rect -1500 436 -1484 464
rect -1456 436 -1440 464
rect -1500 420 -1440 436
rect -1380 464 -1320 480
rect -1380 436 -1364 464
rect -1336 436 -1320 464
rect -1380 420 -1320 436
rect -780 464 -720 480
rect -780 436 -764 464
rect -736 436 -720 464
rect -780 420 -720 436
rect -420 464 -360 480
rect -420 436 -404 464
rect -376 436 -360 464
rect -420 420 -360 436
rect 420 464 480 480
rect 420 436 436 464
rect 464 436 480 464
rect 420 420 480 436
rect 780 464 840 480
rect 780 436 796 464
rect 824 436 840 464
rect 780 420 840 436
rect 1380 464 1440 480
rect 1380 436 1396 464
rect 1424 436 1440 464
rect 1380 420 1440 436
rect 1500 464 1560 480
rect 1500 436 1516 464
rect 1544 436 1560 464
rect 1500 420 1560 436
rect 3420 464 3480 480
rect 3420 436 3436 464
rect 3464 436 3480 464
rect 3420 420 3480 436
rect 3780 464 3840 480
rect 3780 436 3796 464
rect 3824 436 3840 464
rect 3780 420 3840 436
rect -4680 180 -4620 240
rect -3180 224 -3120 240
rect -3180 196 -3164 224
rect -3136 196 -3120 224
rect -3180 180 -3120 196
rect -1020 224 -960 240
rect -1020 196 -1004 224
rect -976 196 -960 224
rect -1020 180 -960 196
rect 1020 224 1080 240
rect 1020 196 1036 224
rect 1064 196 1080 224
rect 1020 180 1080 196
rect 3180 224 3240 240
rect 3180 196 3196 224
rect 3224 196 3240 224
rect 3180 180 3240 196
rect -4680 -300 -4620 0
rect -3300 -6 -3240 0
rect -3300 -294 -3284 -6
rect -3256 -294 -3240 -6
rect -3300 -300 -3240 -294
rect -2820 -6 -2760 0
rect -2820 -294 -2804 -6
rect -2776 -294 -2760 -6
rect -2820 -300 -2760 -294
rect -900 -6 -840 0
rect -900 -294 -884 -6
rect -856 -294 -840 -6
rect -900 -300 -840 -294
rect 900 -6 960 0
rect 900 -294 916 -6
rect 944 -294 960 -6
rect 900 -300 960 -294
rect 2820 -6 2880 0
rect 2820 -294 2836 -6
rect 2864 -294 2880 -6
rect 2820 -300 2880 -294
rect 3300 -6 3360 0
rect 3300 -294 3316 -6
rect 3344 -294 3360 -6
rect 3300 -300 3360 -294
rect -4680 -900 -4620 -600
<< via3 >>
rect -1964 1146 -1936 1434
rect 1996 1146 2024 1434
rect -4004 916 -3976 944
rect -164 916 -136 944
rect 196 916 224 944
rect 4036 916 4064 944
rect -2564 676 -2536 704
rect -2204 676 -2176 704
rect -1604 676 -1576 704
rect 1636 676 1664 704
rect 2236 676 2264 704
rect 2596 676 2624 704
rect -3764 436 -3736 464
rect -3404 436 -3376 464
rect -1364 436 -1336 464
rect -764 436 -736 464
rect -404 436 -376 464
rect 436 436 464 464
rect 796 436 824 464
rect 1396 436 1424 464
rect 3436 436 3464 464
rect 3796 436 3824 464
rect -3164 196 -3136 224
rect -1004 196 -976 224
rect 1036 196 1064 224
rect 3196 196 3224 224
rect -2804 -294 -2776 -6
rect 2836 -294 2864 -6
<< metal4 >>
rect -1980 1434 -1920 1440
rect -1980 1146 -1964 1434
rect -1936 1146 -1920 1434
rect -1980 1140 -1920 1146
rect 1980 1434 2040 1440
rect 1980 1146 1996 1434
rect 2024 1146 2040 1434
rect 1980 1140 2040 1146
rect -4020 944 -3960 960
rect -4020 916 -4004 944
rect -3976 916 -3960 944
rect -4020 900 -3960 916
rect -180 944 -120 960
rect -180 916 -164 944
rect -136 916 -120 944
rect -180 900 -120 916
rect 180 944 240 960
rect 180 916 196 944
rect 224 916 240 944
rect 180 900 240 916
rect 4020 944 4080 960
rect 4020 916 4036 944
rect 4064 916 4080 944
rect 4020 900 4080 916
rect -2580 704 -2520 720
rect -2580 676 -2564 704
rect -2536 676 -2520 704
rect -2580 660 -2520 676
rect -2220 704 -2160 720
rect -2220 676 -2204 704
rect -2176 676 -2160 704
rect -2220 660 -2160 676
rect -1620 704 -1560 720
rect -1620 676 -1604 704
rect -1576 676 -1560 704
rect -1620 660 -1560 676
rect 1620 704 1680 720
rect 1620 676 1636 704
rect 1664 676 1680 704
rect 1620 660 1680 676
rect 2220 704 2280 720
rect 2220 676 2236 704
rect 2264 676 2280 704
rect 2220 660 2280 676
rect 2580 704 2640 720
rect 2580 676 2596 704
rect 2624 676 2640 704
rect 2580 660 2640 676
rect -3780 464 -3720 480
rect -3780 436 -3764 464
rect -3736 436 -3720 464
rect -3780 420 -3720 436
rect -3420 464 -3360 480
rect -3420 436 -3404 464
rect -3376 436 -3360 464
rect -3420 420 -3360 436
rect -1380 464 -1320 480
rect -1380 436 -1364 464
rect -1336 436 -1320 464
rect -1380 420 -1320 436
rect -780 464 -720 480
rect -780 436 -764 464
rect -736 436 -720 464
rect -780 420 -720 436
rect -420 464 -360 480
rect -420 436 -404 464
rect -376 436 -360 464
rect -420 420 -360 436
rect 420 464 480 480
rect 420 436 436 464
rect 464 436 480 464
rect 420 420 480 436
rect 780 464 840 480
rect 780 436 796 464
rect 824 436 840 464
rect 780 420 840 436
rect 1380 464 1440 480
rect 1380 436 1396 464
rect 1424 436 1440 464
rect 1380 420 1440 436
rect 3420 464 3480 480
rect 3420 436 3436 464
rect 3464 436 3480 464
rect 3420 420 3480 436
rect 3780 464 3840 480
rect 3780 436 3796 464
rect 3824 436 3840 464
rect 3780 420 3840 436
rect -3180 224 -3120 240
rect -3180 196 -3164 224
rect -3136 196 -3120 224
rect -3180 180 -3120 196
rect -1020 224 -960 240
rect -1020 196 -1004 224
rect -976 196 -960 224
rect -1020 180 -960 196
rect 1020 224 1080 240
rect 1020 196 1036 224
rect 1064 196 1080 224
rect 1020 180 1080 196
rect 3180 224 3240 240
rect 3180 196 3196 224
rect 3224 196 3240 224
rect 3180 180 3240 196
rect -2820 -6 -2760 0
rect -2820 -294 -2804 -6
rect -2776 -294 -2760 -6
rect -2820 -300 -2760 -294
rect 2820 -6 2880 0
rect 2820 -294 2836 -6
rect 2864 -294 2880 -6
rect 2820 -300 2880 -294
use manf_cell  manf_cell_0
timestamp 1665184495
transform -1 0 660 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_1
timestamp 1665184495
transform -1 0 60 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_2
timestamp 1665184495
transform -1 0 -540 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_3
timestamp 1665184495
transform -1 0 -1140 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_4
timestamp 1665184495
transform -1 0 -1740 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_5
timestamp 1665184495
transform -1 0 -2340 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_6
timestamp 1665184495
transform -1 0 -2940 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_7
timestamp 1665184495
transform 1 0 3000 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_8
timestamp 1665184495
transform 1 0 2400 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_9
timestamp 1665184495
transform 1 0 1800 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_10
timestamp 1665184495
transform 1 0 1200 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_11
timestamp 1665184495
transform 1 0 600 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_12
timestamp 1665184495
transform 1 0 0 0 1 -240
box -3600 -660 -2940 3300
use manf_cell  manf_cell_13
timestamp 1665184495
transform 1 0 -600 0 1 -240
box -3600 -660 -2940 3300
use manf_edge  manf_edge_0
timestamp 1665184495
transform -1 0 900 0 1 -240
box -3780 -660 -3300 3300
use manf_edge  manf_edge_1
timestamp 1665184495
transform 1 0 -840 0 1 -240
box -3780 -660 -3300 3300
<< labels >>
rlabel metal3 s -4650 690 -4650 690 4 x
rlabel metal3 s -4650 450 -4650 450 4 y
rlabel metal3 s -4680 180 -4620 240 4 ip
port 1 nsew
rlabel metal3 s -4680 900 -4620 960 4 im
port 2 nsew
rlabel metal3 s -4680 1140 -4620 1440 4 op
port 3 nsew
rlabel metal3 s -4680 -300 -4620 0 4 om
port 4 nsew
rlabel metal3 s -4680 2640 -4620 2940 4 vdd
port 5 nsew
rlabel metal3 s -4680 2280 -4620 2340 4 gp
port 6 nsew
rlabel metal3 s -4680 1620 -4620 1680 4 bp
port 7 nsew
rlabel metal3 s -4680 2400 -4620 2460 4 vreg
port 8 nsew
rlabel metal3 s -4680 -900 -4620 -600 4 gnd
port 9 nsew
<< end >>
