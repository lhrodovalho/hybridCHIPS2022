* NGSPICE file created from manfvieru.ext - technology: gf180mcuC

.subckt manfvieru_edge gp vreg im ip xm op xp om x y vdd gnd bp
X0 vreg hi hi bp pmos_3p3 w=1.5u l=0.6u
X1 gnd lo lo gnd nmos_3p3 w=1.8u l=0.6u
X2 vdd hih hih vdd pmos_6p0 w=1.8u l=0.6u
C0 vreg hi 0.11fF
C1 hi bp 0.28fF
C2 om xp 0.98fF
C3 xm op 0.98fF
C4 vdd hih 0.45fF
C5 vreg bp 0.23fF
C6 vreg vdd 0.22fF
C7 vreg gp 1.01fF
C8 vreg gnd 0.44fF
C9 bp gnd 4.35fF
C10 vdd gnd 4.01fF
C11 lo gnd 0.84fF
C12 hi gnd 0.46fF
C13 hih gnd 0.46fF
.ends

.subckt manfvieru_cell inl inr out gp vreg op xm im ip xp om x y vdd gnd bp
X0 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X1 out inl vreg bp pmos_3p3 w=1.5u l=0.6u
X2 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X3 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X4 dr inr out gnd nmos_3p3 w=1.8u l=0.6u
X5 dl inl gnd gnd nmos_3p3 w=1.8u l=0.6u
X6 vreg inr out bp pmos_3p3 w=1.5u l=0.6u
X7 gnd inr dr gnd nmos_3p3 w=1.8u l=0.6u
X8 out inl dl gnd nmos_3p3 w=1.8u l=0.6u
X9 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X10 out inr vreg bp pmos_3p3 w=1.5u l=0.6u
X11 vreg inl out bp pmos_3p3 w=1.5u l=0.6u
C0 inl bp 0.32fF
C1 inl op 0.20fF
C2 op xm 1.35fF
C3 bp out 0.15fF
C4 op out 0.12fF
C5 vreg vdd 1.41fF
C6 vdd gp 0.66fF
C7 vreg gp 1.98fF
C8 om inr 0.18fF
C9 inl inr 0.64fF
C10 om inl 0.18fF
C11 out inr 0.20fF
C12 vreg out 0.78fF
C13 om out 0.12fF
C14 bp inr 0.32fF
C15 vreg bp 0.92fF
C16 op inr 0.20fF
C17 inl out 0.18fF
C18 xp om 1.35fF
C19 out gnd 1.80fF
C20 inr gnd 2.38fF
C21 inl gnd 2.39fF
C22 vreg gnd 0.72fF
C23 gp gnd 1.56fF
C24 bp gnd 6.58fF
C25 vdd gnd 6.08fF
C26 dr gnd 0.18fF
C27 dl gnd 0.18fF
.ends

.subckt manfvieru ip im op om vdd gp bp vreg gnd
Xmanfvieru_edge_0 gp vreg im ip xm op xp om x y vdd gnd bp manfvieru_edge
Xmanfvieru_edge_1 gp vreg im ip xm op xp om x y vdd gnd bp manfvieru_edge
Xmanfvieru_cell_0 im y xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_1 y ip xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_2 xp x x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_30 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_3 x om y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_20 im y xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_31 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_4 y y y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_21 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_32 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_10 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_5 op x y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_22 xp x x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_33 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_11 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_7 ip y xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_6 x xm x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_23 y ip xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_12 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_8 y im xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_24 y y y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_9 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_13 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_25 x om y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_14 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_27 op x y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_26 x xm x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_15 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_16 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_17 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_28 ip y xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_18 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_29 y im xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_19 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
X0 om xp mim_2p0fF c_width=199.2u c_length=7.2u
X1 op xm mim_2p0fF c_width=199.2u c_length=7.2u
C0 vreg op 1.05fF
C1 vreg om 0.16fF
C2 vreg x 0.13fF
C3 xm op 52.48fF
C4 op vdd 4.12fF
C5 xm om 0.66fF
C6 xm x 0.20fF
C7 op im 0.52fF
C8 im om 1.05fF
C9 im x 0.15fF
C10 xm ip 1.12fF
C11 op y 1.33fF
C12 y om 1.64fF
C13 x y 0.53fF
C14 op xp 0.67fF
C15 im ip 3.37fF
C16 xp om 52.23fF
C17 x xp 0.29fF
C18 y ip 0.20fF
C19 xp bp 0.11fF
C20 vreg xm 1.31fF
C21 gp op 0.65fF
C22 vreg vdd 0.78fF
C23 ip xp 1.04fF
C24 vreg y 0.20fF
C25 xm vdd 5.42fF
C26 xm im 0.11fF
C27 vreg xp 0.14fF
C28 op om 0.43fF
C29 op x 0.28fF
C30 xm y 0.36fF
C31 op bp 0.13fF
C32 x om 0.41fF
C33 gp vreg -2.47fF
C34 im y 0.15fF
C35 xm xp 0.52fF
C36 op ip 0.71fF
C37 ip om 0.66fF
C38 x ip 0.37fF
C39 im xp 2.13fF
C40 gp xm 0.72fF
C41 gp vdd 0.27fF
C42 y xp 0.72fF
C43 bp gnd 207.63fF
C44 vdd gnd 183.59fF
C45 om gnd 71.62fF
C46 xp gnd 41.51fF
C47 ip gnd 52.08fF
C48 y gnd 63.08fF
C49 x gnd 49.40fF
C50 im gnd 52.06fF
C51 op gnd 56.87fF
C52 xm gnd 35.92fF
C53 vreg gnd 9.16fF
C54 gp gnd 47.13fF
.ends

