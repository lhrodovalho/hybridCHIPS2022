magic
tech gf180mcuC
timestamp 1663179863
<< nwell >>
rect -738 522 -660 642
rect -738 366 -660 498
<< nmos >>
rect -696 -108 -684 -72
<< pmos >>
rect -696 420 -684 450
<< mvpmos >>
rect -696 576 -684 612
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
<< pdiff >>
rect -708 441 -696 450
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 429 -696 435
rect -708 423 -705 429
rect -699 423 -696 429
rect -708 420 -696 423
rect -684 441 -672 450
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 429 -672 435
rect -684 423 -681 429
rect -675 423 -672 429
rect -684 420 -672 423
<< mvpdiff >>
rect -708 609 -696 612
rect -708 603 -705 609
rect -699 603 -696 609
rect -708 597 -696 603
rect -708 591 -705 597
rect -699 591 -696 597
rect -708 585 -696 591
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 576 -696 579
rect -684 609 -672 612
rect -684 603 -681 609
rect -675 603 -672 609
rect -684 597 -672 603
rect -684 591 -681 597
rect -675 591 -672 597
rect -684 585 -672 591
rect -684 579 -681 585
rect -675 579 -672 585
rect -684 576 -672 579
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
<< pdiffc >>
rect -705 435 -699 441
rect -705 423 -699 429
rect -681 435 -675 441
rect -681 423 -675 429
<< mvpdiffc >>
rect -705 603 -699 609
rect -705 591 -699 597
rect -705 579 -699 585
rect -681 603 -675 609
rect -681 591 -675 597
rect -681 579 -675 585
<< psubdiff >>
rect -756 657 -660 660
rect -756 651 -753 657
rect -747 651 -741 657
rect -735 651 -729 657
rect -723 651 -717 657
rect -711 651 -705 657
rect -699 651 -693 657
rect -687 651 -681 657
rect -675 651 -669 657
rect -663 651 -660 657
rect -756 648 -660 651
rect -756 645 -744 648
rect -756 639 -753 645
rect -747 639 -744 645
rect -756 633 -744 639
rect -756 627 -753 633
rect -747 627 -744 633
rect -756 621 -744 627
rect -756 615 -753 621
rect -747 615 -744 621
rect -756 609 -744 615
rect -756 603 -753 609
rect -747 603 -744 609
rect -756 597 -744 603
rect -756 591 -753 597
rect -747 591 -744 597
rect -756 585 -744 591
rect -756 579 -753 585
rect -747 579 -744 585
rect -756 573 -744 579
rect -756 567 -753 573
rect -747 567 -744 573
rect -756 561 -744 567
rect -756 555 -753 561
rect -747 555 -744 561
rect -756 549 -744 555
rect -756 543 -753 549
rect -747 543 -744 549
rect -756 537 -744 543
rect -756 531 -753 537
rect -747 531 -744 537
rect -756 525 -744 531
rect -756 519 -753 525
rect -747 519 -744 525
rect -756 516 -744 519
rect -756 513 -660 516
rect -756 507 -753 513
rect -747 507 -741 513
rect -735 507 -729 513
rect -723 507 -717 513
rect -711 507 -705 513
rect -699 507 -693 513
rect -687 507 -681 513
rect -675 507 -669 513
rect -663 507 -660 513
rect -756 504 -660 507
rect -756 501 -744 504
rect -756 495 -753 501
rect -747 495 -744 501
rect -756 489 -744 495
rect -756 483 -753 489
rect -747 483 -744 489
rect -756 477 -744 483
rect -756 471 -753 477
rect -747 471 -744 477
rect -756 465 -744 471
rect -756 459 -753 465
rect -747 459 -744 465
rect -756 453 -744 459
rect -756 447 -753 453
rect -747 447 -744 453
rect -756 441 -744 447
rect -756 435 -753 441
rect -747 435 -744 441
rect -756 429 -744 435
rect -756 423 -753 429
rect -747 423 -744 429
rect -756 417 -744 423
rect -756 411 -753 417
rect -747 411 -744 417
rect -756 405 -744 411
rect -756 399 -753 405
rect -747 399 -744 405
rect -756 393 -744 399
rect -756 387 -753 393
rect -747 387 -744 393
rect -756 381 -744 387
rect -756 375 -753 381
rect -747 375 -744 381
rect -756 369 -744 375
rect -756 363 -753 369
rect -747 363 -744 369
rect -756 360 -744 363
rect -756 357 -660 360
rect -756 351 -753 357
rect -747 351 -741 357
rect -735 351 -729 357
rect -723 351 -717 357
rect -711 351 -705 357
rect -699 351 -693 357
rect -687 351 -681 357
rect -675 351 -669 357
rect -663 351 -660 357
rect -756 348 -660 351
rect -756 345 -744 348
rect -756 339 -753 345
rect -747 339 -744 345
rect -756 333 -744 339
rect -756 327 -753 333
rect -747 327 -744 333
rect -756 321 -744 327
rect -756 315 -753 321
rect -747 315 -744 321
rect -756 309 -744 315
rect -756 303 -753 309
rect -747 303 -744 309
rect -756 297 -744 303
rect -756 291 -753 297
rect -747 291 -744 297
rect -756 285 -744 291
rect -756 279 -753 285
rect -747 279 -744 285
rect -756 273 -744 279
rect -756 267 -753 273
rect -747 267 -744 273
rect -756 264 -744 267
rect -756 261 -660 264
rect -756 255 -753 261
rect -747 255 -741 261
rect -735 255 -729 261
rect -723 255 -717 261
rect -711 255 -705 261
rect -699 255 -693 261
rect -687 255 -681 261
rect -675 255 -669 261
rect -663 255 -660 261
rect -756 252 -660 255
rect -756 249 -744 252
rect -756 243 -753 249
rect -747 243 -744 249
rect -756 237 -744 243
rect -756 231 -753 237
rect -747 231 -744 237
rect -756 225 -744 231
rect -756 219 -753 225
rect -747 219 -744 225
rect -756 216 -744 219
rect -756 213 -660 216
rect -756 207 -753 213
rect -747 207 -741 213
rect -735 207 -729 213
rect -723 207 -717 213
rect -711 207 -705 213
rect -699 207 -693 213
rect -687 207 -681 213
rect -675 207 -669 213
rect -663 207 -660 213
rect -756 204 -660 207
rect -756 201 -744 204
rect -756 195 -753 201
rect -747 195 -744 201
rect -756 189 -744 195
rect -756 183 -753 189
rect -747 183 -744 189
rect -756 177 -744 183
rect -756 171 -753 177
rect -747 171 -744 177
rect -756 168 -744 171
rect -756 165 -660 168
rect -756 159 -753 165
rect -747 159 -741 165
rect -735 159 -729 165
rect -723 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -660 165
rect -756 156 -660 159
rect -756 153 -744 156
rect -756 147 -753 153
rect -747 147 -744 153
rect -756 141 -744 147
rect -756 135 -753 141
rect -747 135 -744 141
rect -756 129 -744 135
rect -756 123 -753 129
rect -747 123 -744 129
rect -756 120 -744 123
rect -756 117 -660 120
rect -756 111 -753 117
rect -747 111 -741 117
rect -735 111 -729 117
rect -723 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -660 117
rect -756 108 -660 111
rect -756 105 -744 108
rect -756 99 -753 105
rect -747 99 -744 105
rect -756 93 -744 99
rect -756 87 -753 93
rect -747 87 -744 93
rect -756 81 -744 87
rect -756 75 -753 81
rect -747 75 -744 81
rect -756 72 -744 75
rect -756 69 -660 72
rect -756 63 -753 69
rect -747 63 -741 69
rect -735 63 -729 69
rect -723 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -660 69
rect -756 60 -660 63
rect -756 57 -744 60
rect -756 51 -753 57
rect -747 51 -744 57
rect -756 45 -744 51
rect -756 39 -753 45
rect -747 39 -744 45
rect -756 33 -744 39
rect -756 27 -753 33
rect -747 27 -744 33
rect -756 21 -744 27
rect -756 15 -753 21
rect -747 15 -744 21
rect -756 9 -744 15
rect -756 3 -753 9
rect -747 3 -744 9
rect -756 -3 -744 3
rect -756 -9 -753 -3
rect -747 -9 -744 -3
rect -756 -15 -744 -9
rect -756 -21 -753 -15
rect -747 -21 -744 -15
rect -756 -24 -744 -21
rect -756 -27 -660 -24
rect -756 -33 -753 -27
rect -747 -33 -741 -27
rect -735 -33 -729 -27
rect -723 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -39 -744 -36
rect -756 -45 -753 -39
rect -747 -45 -744 -39
rect -756 -51 -744 -45
rect -756 -57 -753 -51
rect -747 -57 -744 -51
rect -756 -63 -744 -57
rect -756 -69 -753 -63
rect -747 -69 -744 -63
rect -756 -75 -744 -69
rect -756 -81 -753 -75
rect -747 -81 -744 -75
rect -756 -87 -744 -81
rect -756 -93 -753 -87
rect -747 -93 -744 -87
rect -756 -99 -744 -93
rect -756 -105 -753 -99
rect -747 -105 -744 -99
rect -756 -111 -744 -105
rect -756 -117 -753 -111
rect -747 -117 -744 -111
rect -756 -120 -744 -117
rect -756 -123 -660 -120
rect -756 -129 -753 -123
rect -747 -129 -741 -123
rect -735 -129 -729 -123
rect -723 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -660 -123
rect -756 -132 -660 -129
<< nsubdiff >>
rect -732 489 -672 492
rect -732 483 -729 489
rect -723 483 -717 489
rect -711 483 -705 489
rect -699 483 -693 489
rect -687 483 -681 489
rect -675 483 -672 489
rect -732 480 -672 483
rect -732 477 -720 480
rect -732 471 -729 477
rect -723 471 -720 477
rect -732 465 -720 471
rect -732 459 -729 465
rect -723 459 -720 465
rect -732 453 -720 459
rect -732 447 -729 453
rect -723 447 -720 453
rect -732 441 -720 447
rect -732 435 -729 441
rect -723 435 -720 441
rect -732 429 -720 435
rect -732 423 -729 429
rect -723 423 -720 429
rect -732 417 -720 423
rect -732 411 -729 417
rect -723 411 -720 417
rect -732 405 -720 411
rect -732 399 -729 405
rect -723 399 -720 405
rect -732 393 -720 399
rect -732 387 -729 393
rect -723 387 -720 393
rect -732 384 -720 387
rect -732 381 -672 384
rect -732 375 -729 381
rect -723 375 -717 381
rect -711 375 -705 381
rect -699 375 -693 381
rect -687 375 -681 381
rect -675 375 -672 381
rect -732 372 -672 375
<< mvnsubdiff >>
rect -732 633 -672 636
rect -732 627 -729 633
rect -723 627 -717 633
rect -711 627 -705 633
rect -699 627 -693 633
rect -687 627 -681 633
rect -675 627 -672 633
rect -732 624 -672 627
rect -732 621 -720 624
rect -732 615 -729 621
rect -723 615 -720 621
rect -732 609 -720 615
rect -732 603 -729 609
rect -723 603 -720 609
rect -732 597 -720 603
rect -732 591 -729 597
rect -723 591 -720 597
rect -732 585 -720 591
rect -732 579 -729 585
rect -723 579 -720 585
rect -732 573 -720 579
rect -732 567 -729 573
rect -723 567 -720 573
rect -732 561 -720 567
rect -732 555 -729 561
rect -723 555 -720 561
rect -732 549 -720 555
rect -732 543 -729 549
rect -723 543 -720 549
rect -732 540 -720 543
rect -732 537 -672 540
rect -732 531 -729 537
rect -723 531 -717 537
rect -711 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -672 537
rect -732 528 -672 531
<< psubdiffcont >>
rect -753 651 -747 657
rect -741 651 -735 657
rect -729 651 -723 657
rect -717 651 -711 657
rect -705 651 -699 657
rect -693 651 -687 657
rect -681 651 -675 657
rect -669 651 -663 657
rect -753 639 -747 645
rect -753 627 -747 633
rect -753 615 -747 621
rect -753 603 -747 609
rect -753 591 -747 597
rect -753 579 -747 585
rect -753 567 -747 573
rect -753 555 -747 561
rect -753 543 -747 549
rect -753 531 -747 537
rect -753 519 -747 525
rect -753 507 -747 513
rect -741 507 -735 513
rect -729 507 -723 513
rect -717 507 -711 513
rect -705 507 -699 513
rect -693 507 -687 513
rect -681 507 -675 513
rect -669 507 -663 513
rect -753 495 -747 501
rect -753 483 -747 489
rect -753 471 -747 477
rect -753 459 -747 465
rect -753 447 -747 453
rect -753 435 -747 441
rect -753 423 -747 429
rect -753 411 -747 417
rect -753 399 -747 405
rect -753 387 -747 393
rect -753 375 -747 381
rect -753 363 -747 369
rect -753 351 -747 357
rect -741 351 -735 357
rect -729 351 -723 357
rect -717 351 -711 357
rect -705 351 -699 357
rect -693 351 -687 357
rect -681 351 -675 357
rect -669 351 -663 357
rect -753 339 -747 345
rect -753 327 -747 333
rect -753 315 -747 321
rect -753 303 -747 309
rect -753 291 -747 297
rect -753 279 -747 285
rect -753 267 -747 273
rect -753 255 -747 261
rect -741 255 -735 261
rect -729 255 -723 261
rect -717 255 -711 261
rect -705 255 -699 261
rect -693 255 -687 261
rect -681 255 -675 261
rect -669 255 -663 261
rect -753 243 -747 249
rect -753 231 -747 237
rect -753 219 -747 225
rect -753 207 -747 213
rect -741 207 -735 213
rect -729 207 -723 213
rect -717 207 -711 213
rect -705 207 -699 213
rect -693 207 -687 213
rect -681 207 -675 213
rect -669 207 -663 213
rect -753 195 -747 201
rect -753 183 -747 189
rect -753 171 -747 177
rect -753 159 -747 165
rect -741 159 -735 165
rect -729 159 -723 165
rect -717 159 -711 165
rect -705 159 -699 165
rect -693 159 -687 165
rect -681 159 -675 165
rect -669 159 -663 165
rect -753 147 -747 153
rect -753 135 -747 141
rect -753 123 -747 129
rect -753 111 -747 117
rect -741 111 -735 117
rect -729 111 -723 117
rect -717 111 -711 117
rect -705 111 -699 117
rect -693 111 -687 117
rect -681 111 -675 117
rect -669 111 -663 117
rect -753 99 -747 105
rect -753 87 -747 93
rect -753 75 -747 81
rect -753 63 -747 69
rect -741 63 -735 69
rect -729 63 -723 69
rect -717 63 -711 69
rect -705 63 -699 69
rect -693 63 -687 69
rect -681 63 -675 69
rect -669 63 -663 69
rect -753 51 -747 57
rect -753 39 -747 45
rect -753 27 -747 33
rect -753 15 -747 21
rect -753 3 -747 9
rect -753 -9 -747 -3
rect -753 -21 -747 -15
rect -753 -33 -747 -27
rect -741 -33 -735 -27
rect -729 -33 -723 -27
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -753 -45 -747 -39
rect -753 -57 -747 -51
rect -753 -69 -747 -63
rect -753 -81 -747 -75
rect -753 -93 -747 -87
rect -753 -105 -747 -99
rect -753 -117 -747 -111
rect -753 -129 -747 -123
rect -741 -129 -735 -123
rect -729 -129 -723 -123
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
<< nsubdiffcont >>
rect -729 483 -723 489
rect -717 483 -711 489
rect -705 483 -699 489
rect -693 483 -687 489
rect -681 483 -675 489
rect -729 471 -723 477
rect -729 459 -723 465
rect -729 447 -723 453
rect -729 435 -723 441
rect -729 423 -723 429
rect -729 411 -723 417
rect -729 399 -723 405
rect -729 387 -723 393
rect -729 375 -723 381
rect -717 375 -711 381
rect -705 375 -699 381
rect -693 375 -687 381
rect -681 375 -675 381
<< mvnsubdiffcont >>
rect -729 627 -723 633
rect -717 627 -711 633
rect -705 627 -699 633
rect -693 627 -687 633
rect -681 627 -675 633
rect -729 615 -723 621
rect -729 603 -723 609
rect -729 591 -723 597
rect -729 579 -723 585
rect -729 567 -723 573
rect -729 555 -723 561
rect -729 543 -723 549
rect -729 531 -723 537
rect -717 531 -711 537
rect -705 531 -699 537
rect -693 531 -687 537
rect -681 531 -675 537
<< polysilicon >>
rect -696 612 -684 618
rect -696 561 -684 576
rect -696 555 -693 561
rect -687 555 -684 561
rect -696 552 -684 555
rect -696 450 -684 456
rect -696 405 -684 420
rect -696 399 -693 405
rect -687 399 -684 405
rect -696 396 -684 399
rect -696 -51 -684 -48
rect -696 -57 -693 -51
rect -687 -57 -684 -51
rect -696 -72 -684 -57
rect -696 -114 -684 -108
<< polycontact >>
rect -693 555 -687 561
rect -693 399 -687 405
rect -693 -57 -687 -51
<< metal1 >>
rect -756 657 -660 660
rect -756 651 -753 657
rect -747 651 -741 657
rect -735 651 -729 657
rect -723 651 -717 657
rect -711 651 -705 657
rect -699 651 -693 657
rect -687 651 -681 657
rect -675 651 -669 657
rect -663 651 -660 657
rect -756 648 -660 651
rect -756 645 -744 648
rect -756 639 -753 645
rect -747 639 -744 645
rect -756 633 -744 639
rect -756 627 -753 633
rect -747 627 -744 633
rect -756 621 -744 627
rect -756 615 -753 621
rect -747 615 -744 621
rect -756 609 -744 615
rect -756 603 -753 609
rect -747 603 -744 609
rect -756 597 -744 603
rect -756 591 -753 597
rect -747 591 -744 597
rect -756 585 -744 591
rect -756 579 -753 585
rect -747 579 -744 585
rect -756 573 -744 579
rect -756 567 -753 573
rect -747 567 -744 573
rect -756 561 -744 567
rect -756 555 -753 561
rect -747 555 -744 561
rect -756 549 -744 555
rect -756 543 -753 549
rect -747 543 -744 549
rect -756 537 -744 543
rect -756 531 -753 537
rect -747 531 -744 537
rect -756 525 -744 531
rect -732 633 -660 636
rect -732 627 -729 633
rect -723 627 -717 633
rect -711 627 -705 633
rect -699 627 -693 633
rect -687 627 -681 633
rect -675 627 -660 633
rect -732 624 -660 627
rect -732 621 -720 624
rect -732 615 -729 621
rect -723 615 -720 621
rect -732 609 -720 615
rect -732 603 -729 609
rect -723 603 -720 609
rect -732 597 -720 603
rect -732 591 -729 597
rect -723 591 -720 597
rect -732 585 -720 591
rect -732 579 -729 585
rect -723 579 -720 585
rect -732 573 -720 579
rect -732 567 -729 573
rect -723 567 -720 573
rect -732 561 -720 567
rect -732 555 -729 561
rect -723 555 -720 561
rect -732 549 -720 555
rect -708 609 -696 612
rect -708 603 -705 609
rect -699 603 -696 609
rect -708 597 -696 603
rect -708 591 -705 597
rect -699 591 -696 597
rect -708 585 -696 591
rect -708 579 -705 585
rect -699 579 -696 585
rect -708 564 -696 579
rect -684 609 -672 612
rect -684 603 -681 609
rect -675 603 -672 609
rect -684 597 -672 603
rect -684 591 -681 597
rect -675 591 -672 597
rect -684 585 -672 591
rect -684 579 -681 585
rect -675 579 -672 585
rect -684 576 -672 579
rect -708 561 -684 564
rect -708 555 -693 561
rect -687 555 -684 561
rect -708 552 -684 555
rect -732 543 -729 549
rect -723 543 -720 549
rect -732 540 -720 543
rect -732 537 -660 540
rect -732 531 -729 537
rect -723 531 -717 537
rect -711 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -660 537
rect -732 528 -660 531
rect -756 519 -753 525
rect -747 519 -744 525
rect -756 516 -744 519
rect -756 513 -660 516
rect -756 507 -753 513
rect -747 507 -741 513
rect -735 507 -729 513
rect -723 507 -717 513
rect -711 507 -705 513
rect -699 507 -693 513
rect -687 507 -681 513
rect -675 507 -669 513
rect -663 507 -660 513
rect -756 504 -660 507
rect -756 501 -744 504
rect -756 495 -753 501
rect -747 495 -744 501
rect -756 489 -744 495
rect -756 483 -753 489
rect -747 483 -744 489
rect -756 477 -744 483
rect -756 471 -753 477
rect -747 471 -744 477
rect -756 465 -744 471
rect -756 459 -753 465
rect -747 459 -744 465
rect -756 453 -744 459
rect -756 447 -753 453
rect -747 447 -744 453
rect -756 441 -744 447
rect -756 435 -753 441
rect -747 435 -744 441
rect -756 429 -744 435
rect -756 423 -753 429
rect -747 423 -744 429
rect -756 417 -744 423
rect -756 411 -753 417
rect -747 411 -744 417
rect -756 405 -744 411
rect -756 399 -753 405
rect -747 399 -744 405
rect -756 393 -744 399
rect -756 387 -753 393
rect -747 387 -744 393
rect -756 381 -744 387
rect -756 375 -753 381
rect -747 375 -744 381
rect -756 369 -744 375
rect -732 489 -672 492
rect -732 483 -729 489
rect -723 483 -717 489
rect -711 483 -705 489
rect -699 483 -693 489
rect -687 483 -681 489
rect -675 483 -672 489
rect -732 480 -672 483
rect -732 477 -720 480
rect -732 471 -729 477
rect -723 471 -720 477
rect -732 465 -720 471
rect -732 459 -729 465
rect -723 459 -720 465
rect -732 453 -720 459
rect -732 447 -729 453
rect -723 447 -720 453
rect -732 441 -720 447
rect -732 435 -729 441
rect -723 435 -720 441
rect -732 429 -720 435
rect -732 423 -729 429
rect -723 423 -720 429
rect -732 417 -720 423
rect -732 411 -729 417
rect -723 411 -720 417
rect -732 405 -720 411
rect -732 399 -729 405
rect -723 399 -720 405
rect -732 393 -720 399
rect -708 441 -696 450
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 429 -696 435
rect -708 423 -705 429
rect -699 423 -696 429
rect -708 408 -696 423
rect -684 441 -672 450
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 429 -672 435
rect -684 423 -681 429
rect -675 423 -672 429
rect -684 420 -672 423
rect -708 405 -684 408
rect -708 399 -693 405
rect -687 399 -684 405
rect -708 396 -684 399
rect -732 387 -729 393
rect -723 387 -720 393
rect -732 384 -720 387
rect -732 381 -660 384
rect -732 375 -729 381
rect -723 375 -717 381
rect -711 375 -705 381
rect -699 375 -693 381
rect -687 375 -681 381
rect -675 375 -660 381
rect -732 372 -660 375
rect -756 363 -753 369
rect -747 363 -744 369
rect -756 360 -744 363
rect -756 357 -660 360
rect -756 351 -753 357
rect -747 351 -741 357
rect -735 351 -729 357
rect -723 351 -717 357
rect -711 351 -705 357
rect -699 351 -693 357
rect -687 351 -681 357
rect -675 351 -669 357
rect -663 351 -660 357
rect -756 348 -660 351
rect -756 345 -744 348
rect -756 339 -753 345
rect -747 339 -744 345
rect -756 333 -744 339
rect -756 327 -753 333
rect -747 327 -744 333
rect -756 321 -744 327
rect -756 315 -753 321
rect -747 315 -744 321
rect -756 309 -744 315
rect -756 303 -753 309
rect -747 303 -744 309
rect -756 297 -744 303
rect -756 291 -753 297
rect -747 291 -744 297
rect -756 285 -744 291
rect -756 279 -753 285
rect -747 279 -744 285
rect -756 273 -744 279
rect -756 267 -753 273
rect -747 267 -744 273
rect -756 264 -744 267
rect -756 261 -660 264
rect -756 255 -753 261
rect -747 255 -741 261
rect -735 255 -729 261
rect -723 255 -717 261
rect -711 255 -705 261
rect -699 255 -693 261
rect -687 255 -681 261
rect -675 255 -669 261
rect -663 255 -660 261
rect -756 252 -660 255
rect -756 249 -744 252
rect -756 243 -753 249
rect -747 243 -744 249
rect -756 237 -744 243
rect -756 231 -753 237
rect -747 231 -744 237
rect -756 225 -744 231
rect -756 219 -753 225
rect -747 219 -744 225
rect -756 216 -744 219
rect -756 213 -660 216
rect -756 207 -753 213
rect -747 207 -741 213
rect -735 207 -729 213
rect -723 207 -717 213
rect -711 207 -705 213
rect -699 207 -693 213
rect -687 207 -681 213
rect -675 207 -669 213
rect -663 207 -660 213
rect -756 204 -660 207
rect -756 201 -744 204
rect -756 195 -753 201
rect -747 195 -744 201
rect -756 189 -744 195
rect -756 183 -753 189
rect -747 183 -744 189
rect -756 177 -744 183
rect -756 171 -753 177
rect -747 171 -744 177
rect -756 168 -744 171
rect -756 165 -660 168
rect -756 159 -753 165
rect -747 159 -741 165
rect -735 159 -729 165
rect -723 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -660 165
rect -756 156 -660 159
rect -756 153 -744 156
rect -756 147 -753 153
rect -747 147 -744 153
rect -756 141 -744 147
rect -756 135 -753 141
rect -747 135 -744 141
rect -756 129 -744 135
rect -756 123 -753 129
rect -747 123 -744 129
rect -756 120 -744 123
rect -756 117 -660 120
rect -756 111 -753 117
rect -747 111 -741 117
rect -735 111 -729 117
rect -723 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -660 117
rect -756 108 -660 111
rect -756 105 -744 108
rect -756 99 -753 105
rect -747 99 -744 105
rect -756 93 -744 99
rect -756 87 -753 93
rect -747 87 -744 93
rect -756 81 -744 87
rect -756 75 -753 81
rect -747 75 -744 81
rect -756 72 -744 75
rect -756 69 -660 72
rect -756 63 -753 69
rect -747 63 -741 69
rect -735 63 -729 69
rect -723 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -660 69
rect -756 60 -660 63
rect -756 57 -744 60
rect -756 51 -753 57
rect -747 51 -744 57
rect -756 45 -744 51
rect -756 39 -753 45
rect -747 39 -744 45
rect -756 33 -744 39
rect -756 27 -753 33
rect -747 27 -744 33
rect -756 21 -744 27
rect -756 15 -753 21
rect -747 15 -744 21
rect -756 9 -744 15
rect -756 3 -753 9
rect -747 3 -744 9
rect -756 -3 -744 3
rect -756 -9 -753 -3
rect -747 -9 -744 -3
rect -756 -15 -744 -9
rect -756 -21 -753 -15
rect -747 -21 -744 -15
rect -756 -24 -744 -21
rect -756 -27 -660 -24
rect -756 -33 -753 -27
rect -747 -33 -741 -27
rect -735 -33 -729 -27
rect -723 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -39 -744 -36
rect -756 -45 -753 -39
rect -747 -45 -744 -39
rect -756 -51 -744 -45
rect -756 -57 -753 -51
rect -747 -57 -744 -51
rect -756 -63 -744 -57
rect -756 -69 -753 -63
rect -747 -69 -744 -63
rect -756 -75 -744 -69
rect -756 -81 -753 -75
rect -747 -81 -744 -75
rect -756 -87 -744 -81
rect -756 -93 -753 -87
rect -747 -93 -744 -87
rect -756 -99 -744 -93
rect -756 -105 -753 -99
rect -747 -105 -744 -99
rect -756 -111 -744 -105
rect -708 -51 -684 -48
rect -708 -57 -693 -51
rect -687 -57 -684 -51
rect -708 -60 -684 -57
rect -708 -75 -696 -60
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -756 -117 -753 -111
rect -747 -117 -744 -111
rect -756 -120 -744 -117
rect -756 -123 -660 -120
rect -756 -129 -753 -123
rect -747 -129 -741 -123
rect -735 -129 -729 -123
rect -723 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -660 -123
rect -756 -132 -660 -129
<< via1 >>
rect -681 627 -675 633
rect -681 603 -675 609
rect -681 591 -675 597
rect -681 579 -675 585
rect -681 435 -675 441
rect -681 423 -675 429
rect -729 375 -723 381
rect -681 351 -675 357
rect -681 255 -675 261
rect -681 207 -675 213
rect -681 159 -675 165
rect -681 111 -675 117
rect -681 63 -675 69
rect -681 -33 -675 -27
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -681 -129 -675 -123
<< metal2 >>
rect -684 633 -672 636
rect -684 627 -681 633
rect -675 627 -672 633
rect -684 609 -672 627
rect -684 603 -681 609
rect -675 603 -672 609
rect -684 597 -672 603
rect -684 591 -681 597
rect -675 591 -672 597
rect -684 585 -672 591
rect -684 579 -681 585
rect -675 579 -672 585
rect -684 576 -672 579
rect -708 537 -696 540
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 489 -696 531
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 480 -696 483
rect -684 489 -672 492
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 441 -672 483
rect -684 435 -681 441
rect -675 435 -672 441
rect -684 429 -672 435
rect -684 423 -681 429
rect -675 423 -672 429
rect -684 420 -672 423
rect -732 381 -720 384
rect -732 375 -729 381
rect -723 375 -720 381
rect -732 372 -720 375
rect -684 357 -672 360
rect -684 351 -681 357
rect -675 351 -672 357
rect -684 261 -672 351
rect -684 255 -681 261
rect -675 255 -672 261
rect -684 213 -672 255
rect -684 207 -681 213
rect -675 207 -672 213
rect -684 165 -672 207
rect -684 159 -681 165
rect -675 159 -672 165
rect -684 117 -672 159
rect -684 111 -681 117
rect -675 111 -672 117
rect -684 69 -672 111
rect -684 63 -681 69
rect -675 63 -672 69
rect -684 -27 -672 63
rect -684 -33 -681 -27
rect -675 -33 -672 -27
rect -684 -75 -672 -33
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -123 -672 -105
rect -684 -129 -681 -123
rect -675 -129 -672 -123
rect -684 -132 -672 -129
<< via2 >>
rect -681 627 -675 633
rect -681 603 -675 609
rect -681 591 -675 597
rect -681 579 -675 585
rect -705 531 -699 537
rect -705 483 -699 489
rect -681 483 -675 489
rect -729 375 -723 381
rect -681 351 -675 357
rect -681 255 -675 261
rect -681 207 -675 213
rect -681 159 -675 165
rect -681 111 -675 117
rect -681 63 -675 69
rect -681 -33 -675 -27
rect -681 -129 -675 -123
<< metal3 >>
rect -756 633 -660 636
rect -756 627 -681 633
rect -675 627 -660 633
rect -756 609 -660 627
rect -756 603 -681 609
rect -675 603 -660 609
rect -756 597 -660 603
rect -756 591 -681 597
rect -675 591 -660 597
rect -756 585 -660 591
rect -756 579 -681 585
rect -675 579 -660 585
rect -756 576 -660 579
rect -756 537 -660 540
rect -756 531 -705 537
rect -699 531 -660 537
rect -756 522 -660 531
rect -756 504 -660 516
rect -756 489 -660 498
rect -756 483 -705 489
rect -699 483 -681 489
rect -675 483 -660 489
rect -756 480 -660 483
rect -756 381 -660 384
rect -756 375 -729 381
rect -723 375 -660 381
rect -756 372 -660 375
rect -756 357 -660 360
rect -756 351 -681 357
rect -675 351 -660 357
rect -756 348 -660 351
rect -756 276 -660 336
rect -756 261 -660 264
rect -756 255 -681 261
rect -675 255 -660 261
rect -756 252 -660 255
rect -756 228 -660 240
rect -756 213 -660 216
rect -756 207 -681 213
rect -675 207 -660 213
rect -756 204 -660 207
rect -756 180 -660 192
rect -756 165 -660 168
rect -756 159 -681 165
rect -675 159 -660 165
rect -756 156 -660 159
rect -756 132 -660 144
rect -756 117 -660 120
rect -756 111 -681 117
rect -675 111 -660 117
rect -756 108 -660 111
rect -756 84 -660 96
rect -756 69 -660 72
rect -756 63 -681 69
rect -675 63 -660 69
rect -756 60 -660 63
rect -756 -12 -660 48
rect -756 -27 -660 -24
rect -756 -33 -681 -27
rect -675 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -123 -660 -72
rect -756 -129 -681 -123
rect -675 -129 -660 -123
rect -756 -132 -660 -129
<< labels >>
rlabel metal3 -756 576 -660 636 0 vdd
port 1 nsew
rlabel metal3 -756 528 -660 540 0 vreg
port 2 nsew
rlabel metal3 -756 504 -660 516 0 gp
port 3 nsew
rlabel metal3 -756 372 -660 384 0 bp
port 4 nsew
rlabel metal3 -756 276 -660 336 0 op
port 5 nsew
rlabel metal3 -756 228 -660 240 0 im
port 6 nsew
rlabel metal3 -756 180 -660 192 0 x
port 7 nsew
rlabel metal3 -756 132 -660 144 0 y
port 8 nsew
rlabel metal3 -756 84 -660 96 0 ip
port 9 nsew
rlabel metal3 -756 -12 -660 48 0 om
port 10 nsew
rlabel metal3 -756 -132 -660 -72 0 gnd
port 11 nsew
rlabel metal1 -708 552 -696 564 1 hih
rlabel metal1 -708 396 -696 408 0 hi
rlabel metal1 -708 -60 -696 -48 0 lo
<< end >>
