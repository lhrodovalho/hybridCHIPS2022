magic
tech gf180mcuC
timestamp 1663277574
<< nwell >>
rect -720 426 -588 546
rect -720 270 -588 402
<< nmos >>
rect -696 -108 -684 -72
rect -672 -108 -660 -72
rect -648 -108 -636 -72
rect -624 -108 -612 -72
<< pmos >>
rect -696 324 -684 354
rect -672 324 -660 354
rect -648 324 -636 354
rect -624 324 -612 354
<< mvpmos >>
rect -696 480 -684 516
rect -672 480 -660 516
rect -648 480 -636 516
rect -624 480 -612 516
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
<< pdiff >>
rect -708 345 -696 354
rect -708 339 -705 345
rect -699 339 -696 345
rect -708 333 -696 339
rect -708 327 -705 333
rect -699 327 -696 333
rect -708 324 -696 327
rect -684 345 -672 354
rect -684 339 -681 345
rect -675 339 -672 345
rect -684 333 -672 339
rect -684 327 -681 333
rect -675 327 -672 333
rect -684 324 -672 327
rect -660 345 -648 354
rect -660 339 -657 345
rect -651 339 -648 345
rect -660 333 -648 339
rect -660 327 -657 333
rect -651 327 -648 333
rect -660 324 -648 327
rect -636 345 -624 354
rect -636 339 -633 345
rect -627 339 -624 345
rect -636 333 -624 339
rect -636 327 -633 333
rect -627 327 -624 333
rect -636 324 -624 327
rect -612 345 -600 354
rect -612 339 -609 345
rect -603 339 -600 345
rect -612 333 -600 339
rect -612 327 -609 333
rect -603 327 -600 333
rect -612 324 -600 327
<< mvpdiff >>
rect -708 513 -696 516
rect -708 507 -705 513
rect -699 507 -696 513
rect -708 501 -696 507
rect -708 495 -705 501
rect -699 495 -696 501
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 480 -696 483
rect -684 513 -672 516
rect -684 507 -681 513
rect -675 507 -672 513
rect -684 501 -672 507
rect -684 495 -681 501
rect -675 495 -672 501
rect -684 489 -672 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -660 513 -648 516
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 501 -648 507
rect -660 495 -657 501
rect -651 495 -648 501
rect -660 489 -648 495
rect -660 483 -657 489
rect -651 483 -648 489
rect -660 480 -648 483
rect -636 513 -624 516
rect -636 507 -633 513
rect -627 507 -624 513
rect -636 501 -624 507
rect -636 495 -633 501
rect -627 495 -624 501
rect -636 489 -624 495
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 480 -624 483
rect -612 513 -600 516
rect -612 507 -609 513
rect -603 507 -600 513
rect -612 501 -600 507
rect -612 495 -609 501
rect -603 495 -600 501
rect -612 489 -600 495
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 480 -600 483
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -633 -81 -627 -75
rect -633 -93 -627 -87
rect -633 -105 -627 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
<< pdiffc >>
rect -705 339 -699 345
rect -705 327 -699 333
rect -681 339 -675 345
rect -681 327 -675 333
rect -657 339 -651 345
rect -657 327 -651 333
rect -633 339 -627 345
rect -633 327 -627 333
rect -609 339 -603 345
rect -609 327 -603 333
<< mvpdiffc >>
rect -705 507 -699 513
rect -705 495 -699 501
rect -705 483 -699 489
rect -681 507 -675 513
rect -681 495 -675 501
rect -681 483 -675 489
rect -657 507 -651 513
rect -657 495 -651 501
rect -657 483 -651 489
rect -633 507 -627 513
rect -633 495 -627 501
rect -633 483 -627 489
rect -609 507 -603 513
rect -609 495 -603 501
rect -609 483 -603 489
<< psubdiff >>
rect -720 561 -588 564
rect -720 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -657 561
rect -651 555 -645 561
rect -639 555 -633 561
rect -627 555 -621 561
rect -615 555 -609 561
rect -603 555 -597 561
rect -591 555 -588 561
rect -720 552 -588 555
rect -720 417 -588 420
rect -720 411 -717 417
rect -711 411 -705 417
rect -699 411 -693 417
rect -687 411 -681 417
rect -675 411 -669 417
rect -663 411 -657 417
rect -651 411 -645 417
rect -639 411 -633 417
rect -627 411 -621 417
rect -615 411 -609 417
rect -603 411 -597 417
rect -591 411 -588 417
rect -720 408 -588 411
rect -720 261 -588 264
rect -720 255 -717 261
rect -711 255 -705 261
rect -699 255 -693 261
rect -687 255 -681 261
rect -675 255 -669 261
rect -663 255 -657 261
rect -651 255 -645 261
rect -639 255 -633 261
rect -627 255 -621 261
rect -615 255 -609 261
rect -603 255 -597 261
rect -591 255 -588 261
rect -720 252 -588 255
rect -720 165 -588 168
rect -720 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -657 165
rect -651 159 -645 165
rect -639 159 -633 165
rect -627 159 -621 165
rect -615 159 -609 165
rect -603 159 -597 165
rect -591 159 -588 165
rect -720 156 -588 159
rect -720 117 -588 120
rect -720 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -657 117
rect -651 111 -645 117
rect -639 111 -633 117
rect -627 111 -621 117
rect -615 111 -609 117
rect -603 111 -597 117
rect -591 111 -588 117
rect -720 108 -588 111
rect -720 69 -588 72
rect -720 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -657 69
rect -651 63 -645 69
rect -639 63 -633 69
rect -627 63 -621 69
rect -615 63 -609 69
rect -603 63 -597 69
rect -591 63 -588 69
rect -720 60 -588 63
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< nsubdiff >>
rect -708 393 -600 396
rect -708 387 -705 393
rect -699 387 -693 393
rect -687 387 -681 393
rect -675 387 -669 393
rect -663 387 -657 393
rect -651 387 -645 393
rect -639 387 -633 393
rect -627 387 -621 393
rect -615 387 -609 393
rect -603 387 -600 393
rect -708 384 -600 387
rect -708 285 -600 288
rect -708 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -669 285
rect -663 279 -657 285
rect -651 279 -645 285
rect -639 279 -633 285
rect -627 279 -621 285
rect -615 279 -609 285
rect -603 279 -600 285
rect -708 276 -600 279
<< mvnsubdiff >>
rect -708 537 -600 540
rect -708 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -669 537
rect -663 531 -657 537
rect -651 531 -645 537
rect -639 531 -633 537
rect -627 531 -621 537
rect -615 531 -609 537
rect -603 531 -600 537
rect -708 528 -600 531
rect -708 441 -600 444
rect -708 435 -705 441
rect -699 435 -693 441
rect -687 435 -681 441
rect -675 435 -669 441
rect -663 435 -657 441
rect -651 435 -645 441
rect -639 435 -633 441
rect -627 435 -621 441
rect -615 435 -609 441
rect -603 435 -600 441
rect -708 432 -600 435
<< psubdiffcont >>
rect -717 555 -711 561
rect -705 555 -699 561
rect -693 555 -687 561
rect -681 555 -675 561
rect -669 555 -663 561
rect -657 555 -651 561
rect -645 555 -639 561
rect -633 555 -627 561
rect -621 555 -615 561
rect -609 555 -603 561
rect -597 555 -591 561
rect -717 411 -711 417
rect -705 411 -699 417
rect -693 411 -687 417
rect -681 411 -675 417
rect -669 411 -663 417
rect -657 411 -651 417
rect -645 411 -639 417
rect -633 411 -627 417
rect -621 411 -615 417
rect -609 411 -603 417
rect -597 411 -591 417
rect -717 255 -711 261
rect -705 255 -699 261
rect -693 255 -687 261
rect -681 255 -675 261
rect -669 255 -663 261
rect -657 255 -651 261
rect -645 255 -639 261
rect -633 255 -627 261
rect -621 255 -615 261
rect -609 255 -603 261
rect -597 255 -591 261
rect -717 159 -711 165
rect -705 159 -699 165
rect -693 159 -687 165
rect -681 159 -675 165
rect -669 159 -663 165
rect -657 159 -651 165
rect -645 159 -639 165
rect -633 159 -627 165
rect -621 159 -615 165
rect -609 159 -603 165
rect -597 159 -591 165
rect -717 111 -711 117
rect -705 111 -699 117
rect -693 111 -687 117
rect -681 111 -675 117
rect -669 111 -663 117
rect -657 111 -651 117
rect -645 111 -639 117
rect -633 111 -627 117
rect -621 111 -615 117
rect -609 111 -603 117
rect -597 111 -591 117
rect -717 63 -711 69
rect -705 63 -699 69
rect -693 63 -687 69
rect -681 63 -675 69
rect -669 63 -663 69
rect -657 63 -651 69
rect -645 63 -639 69
rect -633 63 -627 69
rect -621 63 -615 69
rect -609 63 -603 69
rect -597 63 -591 69
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -657 -33 -651 -27
rect -645 -33 -639 -27
rect -633 -33 -627 -27
rect -621 -33 -615 -27
rect -609 -33 -603 -27
rect -597 -33 -591 -27
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
rect -657 -129 -651 -123
rect -645 -129 -639 -123
rect -633 -129 -627 -123
rect -621 -129 -615 -123
rect -609 -129 -603 -123
rect -597 -129 -591 -123
<< nsubdiffcont >>
rect -705 387 -699 393
rect -693 387 -687 393
rect -681 387 -675 393
rect -669 387 -663 393
rect -657 387 -651 393
rect -645 387 -639 393
rect -633 387 -627 393
rect -621 387 -615 393
rect -609 387 -603 393
rect -705 279 -699 285
rect -693 279 -687 285
rect -681 279 -675 285
rect -669 279 -663 285
rect -657 279 -651 285
rect -645 279 -639 285
rect -633 279 -627 285
rect -621 279 -615 285
rect -609 279 -603 285
<< mvnsubdiffcont >>
rect -705 531 -699 537
rect -693 531 -687 537
rect -681 531 -675 537
rect -669 531 -663 537
rect -657 531 -651 537
rect -645 531 -639 537
rect -633 531 -627 537
rect -621 531 -615 537
rect -609 531 -603 537
rect -705 435 -699 441
rect -693 435 -687 441
rect -681 435 -675 441
rect -669 435 -663 441
rect -657 435 -651 441
rect -645 435 -639 441
rect -633 435 -627 441
rect -621 435 -615 441
rect -609 435 -603 441
<< polysilicon >>
rect -696 516 -684 522
rect -672 516 -660 522
rect -648 516 -636 522
rect -624 516 -612 522
rect -696 468 -684 480
rect -672 468 -660 480
rect -648 468 -636 480
rect -624 468 -612 480
rect -696 465 -612 468
rect -696 459 -693 465
rect -687 459 -681 465
rect -675 459 -669 465
rect -663 459 -657 465
rect -651 459 -645 465
rect -639 459 -633 465
rect -627 459 -621 465
rect -615 459 -612 465
rect -696 456 -612 459
rect -696 354 -684 360
rect -672 354 -660 360
rect -648 354 -636 360
rect -624 354 -612 360
rect -696 312 -684 324
rect -672 312 -660 324
rect -696 309 -660 312
rect -696 303 -693 309
rect -687 303 -681 309
rect -675 303 -669 309
rect -663 303 -660 309
rect -696 300 -660 303
rect -648 312 -636 324
rect -624 312 -612 324
rect -648 309 -612 312
rect -648 303 -645 309
rect -639 303 -633 309
rect -627 303 -621 309
rect -615 303 -612 309
rect -648 300 -612 303
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -696 -72 -684 -60
rect -672 -72 -660 -60
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -648 -72 -636 -60
rect -624 -72 -612 -60
rect -696 -114 -684 -108
rect -672 -114 -660 -108
rect -648 -114 -636 -108
rect -624 -114 -612 -108
<< polycontact >>
rect -693 459 -687 465
rect -681 459 -675 465
rect -669 459 -663 465
rect -657 459 -651 465
rect -645 459 -639 465
rect -633 459 -627 465
rect -621 459 -615 465
rect -693 303 -687 309
rect -681 303 -675 309
rect -669 303 -663 309
rect -645 303 -639 309
rect -633 303 -627 309
rect -621 303 -615 309
rect -693 -57 -687 -51
rect -681 -57 -675 -51
rect -669 -57 -663 -51
rect -645 -57 -639 -51
rect -633 -57 -627 -51
rect -621 -57 -615 -51
<< metal1 >>
rect -720 561 -588 564
rect -720 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -657 561
rect -651 555 -645 561
rect -639 555 -633 561
rect -627 555 -621 561
rect -615 555 -609 561
rect -603 555 -597 561
rect -591 555 -588 561
rect -720 552 -588 555
rect -720 537 -588 540
rect -720 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -669 537
rect -663 531 -657 537
rect -651 531 -645 537
rect -639 531 -633 537
rect -627 531 -621 537
rect -615 531 -609 537
rect -603 531 -588 537
rect -720 528 -588 531
rect -708 513 -696 516
rect -708 507 -705 513
rect -699 507 -696 513
rect -708 501 -696 507
rect -708 495 -705 501
rect -699 495 -696 501
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 480 -696 483
rect -684 513 -672 516
rect -684 507 -681 513
rect -675 507 -672 513
rect -684 501 -672 507
rect -684 495 -681 501
rect -675 495 -672 501
rect -684 489 -672 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -660 513 -648 516
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 501 -648 507
rect -660 495 -657 501
rect -651 495 -648 501
rect -660 489 -648 495
rect -660 483 -657 489
rect -651 483 -648 489
rect -660 480 -648 483
rect -636 513 -624 516
rect -636 507 -633 513
rect -627 507 -624 513
rect -636 501 -624 507
rect -636 495 -633 501
rect -627 495 -624 501
rect -636 489 -624 495
rect -636 483 -633 489
rect -627 483 -624 489
rect -636 480 -624 483
rect -612 513 -600 516
rect -612 507 -609 513
rect -603 507 -600 513
rect -612 501 -600 507
rect -612 495 -609 501
rect -603 495 -600 501
rect -612 489 -600 495
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 480 -600 483
rect -696 465 -612 468
rect -696 459 -693 465
rect -687 459 -681 465
rect -675 459 -669 465
rect -663 459 -657 465
rect -651 459 -645 465
rect -639 459 -633 465
rect -627 459 -621 465
rect -615 459 -612 465
rect -696 456 -612 459
rect -720 441 -588 444
rect -720 435 -705 441
rect -699 435 -693 441
rect -687 435 -681 441
rect -675 435 -669 441
rect -663 435 -657 441
rect -651 435 -645 441
rect -639 435 -633 441
rect -627 435 -621 441
rect -615 435 -609 441
rect -603 435 -588 441
rect -720 432 -588 435
rect -720 417 -588 420
rect -720 411 -717 417
rect -711 411 -705 417
rect -699 411 -693 417
rect -687 411 -681 417
rect -675 411 -669 417
rect -663 411 -657 417
rect -651 411 -645 417
rect -639 411 -633 417
rect -627 411 -621 417
rect -615 411 -609 417
rect -603 411 -597 417
rect -591 411 -588 417
rect -720 408 -588 411
rect -720 393 -588 396
rect -720 387 -705 393
rect -699 387 -693 393
rect -687 387 -681 393
rect -675 387 -669 393
rect -663 387 -657 393
rect -651 387 -645 393
rect -639 387 -633 393
rect -627 387 -621 393
rect -615 387 -609 393
rect -603 387 -588 393
rect -720 384 -588 387
rect -708 369 -600 372
rect -708 363 -705 369
rect -699 363 -657 369
rect -651 363 -609 369
rect -603 363 -600 369
rect -708 360 -600 363
rect -708 357 -696 360
rect -708 351 -705 357
rect -699 351 -696 357
rect -660 357 -648 360
rect -708 345 -696 351
rect -708 339 -705 345
rect -699 339 -696 345
rect -708 333 -696 339
rect -708 327 -705 333
rect -699 327 -696 333
rect -708 324 -696 327
rect -684 345 -672 354
rect -684 339 -681 345
rect -675 339 -672 345
rect -684 333 -672 339
rect -684 327 -681 333
rect -675 327 -672 333
rect -684 324 -672 327
rect -660 351 -657 357
rect -651 351 -648 357
rect -612 357 -600 360
rect -660 345 -648 351
rect -660 339 -657 345
rect -651 339 -648 345
rect -660 333 -648 339
rect -660 327 -657 333
rect -651 327 -648 333
rect -660 324 -648 327
rect -636 345 -624 354
rect -636 339 -633 345
rect -627 339 -624 345
rect -636 333 -624 339
rect -636 327 -633 333
rect -627 327 -624 333
rect -636 324 -624 327
rect -612 351 -609 357
rect -603 351 -600 357
rect -612 345 -600 351
rect -612 339 -609 345
rect -603 339 -600 345
rect -612 333 -600 339
rect -612 327 -609 333
rect -603 327 -600 333
rect -612 324 -600 327
rect -696 309 -660 312
rect -696 303 -693 309
rect -687 303 -681 309
rect -675 303 -669 309
rect -663 303 -660 309
rect -696 300 -660 303
rect -648 309 -612 312
rect -648 303 -645 309
rect -639 303 -633 309
rect -627 303 -621 309
rect -615 303 -612 309
rect -648 300 -612 303
rect -720 285 -588 288
rect -720 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -669 285
rect -663 279 -657 285
rect -651 279 -645 285
rect -639 279 -633 285
rect -627 279 -621 285
rect -615 279 -609 285
rect -603 279 -588 285
rect -720 276 -588 279
rect -720 261 -588 264
rect -720 255 -717 261
rect -711 255 -705 261
rect -699 255 -693 261
rect -687 255 -681 261
rect -675 255 -669 261
rect -663 255 -657 261
rect -651 255 -645 261
rect -639 255 -633 261
rect -627 255 -621 261
rect -615 255 -609 261
rect -603 255 -597 261
rect -591 255 -588 261
rect -720 252 -588 255
rect -720 165 -588 168
rect -720 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -657 165
rect -651 159 -645 165
rect -639 159 -633 165
rect -627 159 -621 165
rect -615 159 -609 165
rect -603 159 -597 165
rect -591 159 -588 165
rect -720 156 -588 159
rect -720 117 -588 120
rect -720 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -657 117
rect -651 111 -645 117
rect -639 111 -633 117
rect -627 111 -621 117
rect -615 111 -609 117
rect -603 111 -597 117
rect -591 111 -588 117
rect -720 108 -588 111
rect -720 69 -588 72
rect -720 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -657 69
rect -651 63 -645 69
rect -639 63 -633 69
rect -627 63 -621 69
rect -615 63 -609 69
rect -603 63 -597 69
rect -591 63 -588 69
rect -720 60 -588 63
rect -720 -27 -588 -24
rect -720 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -657 -27
rect -651 -33 -645 -27
rect -639 -33 -633 -27
rect -627 -33 -621 -27
rect -615 -33 -609 -27
rect -603 -33 -597 -27
rect -591 -33 -588 -27
rect -720 -36 -588 -33
rect -696 -51 -660 -48
rect -696 -57 -693 -51
rect -687 -57 -681 -51
rect -675 -57 -669 -51
rect -663 -57 -660 -51
rect -696 -60 -660 -57
rect -648 -51 -612 -48
rect -648 -57 -645 -51
rect -639 -57 -633 -51
rect -627 -57 -621 -51
rect -615 -57 -612 -51
rect -648 -60 -612 -57
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -660 -75 -648 -72
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -636 -75 -624 -72
rect -636 -81 -633 -75
rect -627 -81 -624 -75
rect -636 -87 -624 -81
rect -636 -93 -633 -87
rect -627 -93 -624 -87
rect -636 -99 -624 -93
rect -636 -105 -633 -99
rect -627 -105 -624 -99
rect -636 -108 -624 -105
rect -612 -75 -600 -72
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -612 -108 -600 -105
rect -720 -123 -588 -120
rect -720 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -657 -123
rect -651 -129 -645 -123
rect -639 -129 -633 -123
rect -627 -129 -621 -123
rect -615 -129 -609 -123
rect -603 -129 -597 -123
rect -591 -129 -588 -123
rect -720 -132 -588 -129
<< via1 >>
rect -705 531 -699 537
rect -657 531 -651 537
rect -609 531 -603 537
rect -705 507 -699 513
rect -705 495 -699 501
rect -705 483 -699 489
rect -681 507 -675 513
rect -681 495 -675 501
rect -681 483 -675 489
rect -657 507 -651 513
rect -657 495 -651 501
rect -657 483 -651 489
rect -633 507 -627 513
rect -633 495 -627 501
rect -633 483 -627 489
rect -609 507 -603 513
rect -609 495 -603 501
rect -609 483 -603 489
rect -657 459 -651 465
rect -705 363 -699 369
rect -657 363 -651 369
rect -609 363 -603 369
rect -705 351 -699 357
rect -705 339 -699 345
rect -705 327 -699 333
rect -681 339 -675 345
rect -681 327 -675 333
rect -657 351 -651 357
rect -633 339 -627 345
rect -633 327 -627 333
rect -609 351 -603 357
rect -609 339 -603 345
rect -609 327 -603 333
rect -681 303 -675 309
rect -633 303 -627 309
rect -705 279 -699 285
rect -609 279 -603 285
rect -705 255 -699 261
rect -609 255 -603 261
rect -705 159 -699 165
rect -609 159 -603 165
rect -705 111 -699 117
rect -609 111 -603 117
rect -705 63 -699 69
rect -609 63 -603 69
rect -705 -33 -699 -27
rect -609 -33 -603 -27
rect -681 -57 -675 -51
rect -633 -57 -627 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -657 -81 -651 -75
rect -657 -93 -651 -87
rect -657 -105 -651 -99
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal2 >>
rect -708 537 -696 540
rect -708 531 -705 537
rect -699 531 -696 537
rect -708 513 -696 531
rect -660 537 -648 540
rect -660 531 -657 537
rect -651 531 -648 537
rect -708 507 -705 513
rect -699 507 -696 513
rect -708 501 -696 507
rect -708 495 -705 501
rect -699 495 -696 501
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 480 -696 483
rect -684 513 -672 516
rect -684 507 -681 513
rect -675 507 -672 513
rect -684 501 -672 507
rect -684 495 -681 501
rect -675 495 -672 501
rect -684 489 -672 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 441 -672 483
rect -660 513 -648 531
rect -612 537 -600 540
rect -612 531 -609 537
rect -603 531 -600 537
rect -660 507 -657 513
rect -651 507 -648 513
rect -660 501 -648 507
rect -660 495 -657 501
rect -651 495 -648 501
rect -660 489 -648 495
rect -660 483 -657 489
rect -651 483 -648 489
rect -660 480 -648 483
rect -636 513 -624 516
rect -636 507 -633 513
rect -627 507 -624 513
rect -636 501 -624 507
rect -636 495 -633 501
rect -627 495 -624 501
rect -636 489 -624 495
rect -636 483 -633 489
rect -627 483 -624 489
rect -660 465 -648 468
rect -660 459 -657 465
rect -651 459 -648 465
rect -660 456 -648 459
rect -684 435 -681 441
rect -675 435 -672 441
rect -708 393 -696 396
rect -708 387 -705 393
rect -699 387 -696 393
rect -708 369 -696 387
rect -684 393 -672 435
rect -636 441 -624 483
rect -612 513 -600 531
rect -612 507 -609 513
rect -603 507 -600 513
rect -612 501 -600 507
rect -612 495 -609 501
rect -603 495 -600 501
rect -612 489 -600 495
rect -612 483 -609 489
rect -603 483 -600 489
rect -612 480 -600 483
rect -636 435 -633 441
rect -627 435 -624 441
rect -684 387 -681 393
rect -675 387 -672 393
rect -684 384 -672 387
rect -660 393 -648 396
rect -660 387 -657 393
rect -651 387 -648 393
rect -708 363 -705 369
rect -699 363 -696 369
rect -708 357 -696 363
rect -708 351 -705 357
rect -699 351 -696 357
rect -660 369 -648 387
rect -636 393 -624 435
rect -636 387 -633 393
rect -627 387 -624 393
rect -636 384 -624 387
rect -612 393 -600 396
rect -612 387 -609 393
rect -603 387 -600 393
rect -660 363 -657 369
rect -651 363 -648 369
rect -660 357 -648 363
rect -708 345 -696 351
rect -708 339 -705 345
rect -699 339 -696 345
rect -708 333 -696 339
rect -708 327 -705 333
rect -699 327 -696 333
rect -708 324 -696 327
rect -684 345 -672 354
rect -660 351 -657 357
rect -651 351 -648 357
rect -612 369 -600 387
rect -612 363 -609 369
rect -603 363 -600 369
rect -612 357 -600 363
rect -660 348 -648 351
rect -684 339 -681 345
rect -675 339 -672 345
rect -684 336 -672 339
rect -636 345 -624 354
rect -636 339 -633 345
rect -627 339 -624 345
rect -636 336 -624 339
rect -684 333 -624 336
rect -684 327 -681 333
rect -675 327 -633 333
rect -627 327 -624 333
rect -684 324 -624 327
rect -612 351 -609 357
rect -603 351 -600 357
rect -612 345 -600 351
rect -612 339 -609 345
rect -603 339 -600 345
rect -612 333 -600 339
rect -612 327 -609 333
rect -603 327 -600 333
rect -612 324 -600 327
rect -684 309 -672 312
rect -684 303 -681 309
rect -675 303 -672 309
rect -684 300 -672 303
rect -708 285 -696 288
rect -708 279 -705 285
rect -699 279 -696 285
rect -708 276 -696 279
rect -708 261 -696 264
rect -708 255 -705 261
rect -699 255 -696 261
rect -708 165 -696 255
rect -708 159 -705 165
rect -699 159 -696 165
rect -708 117 -696 159
rect -708 111 -705 117
rect -699 111 -696 117
rect -708 69 -696 111
rect -708 63 -705 69
rect -699 63 -696 69
rect -708 -27 -696 63
rect -708 -33 -705 -27
rect -699 -33 -696 -27
rect -708 -75 -696 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -123 -696 -105
rect -660 -75 -648 324
rect -636 309 -624 312
rect -636 303 -633 309
rect -627 303 -624 309
rect -636 300 -624 303
rect -612 285 -600 288
rect -612 279 -609 285
rect -603 279 -600 285
rect -612 276 -600 279
rect -612 261 -600 264
rect -612 255 -609 261
rect -603 255 -600 261
rect -612 165 -600 255
rect -612 159 -609 165
rect -603 159 -600 165
rect -612 117 -600 159
rect -612 111 -609 117
rect -603 111 -600 117
rect -612 69 -600 111
rect -612 63 -609 69
rect -603 63 -600 69
rect -612 -27 -600 63
rect -612 -33 -609 -27
rect -603 -33 -600 -27
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -660 -81 -657 -75
rect -651 -81 -648 -75
rect -660 -87 -648 -81
rect -660 -93 -657 -87
rect -651 -93 -648 -87
rect -660 -99 -648 -93
rect -660 -105 -657 -99
rect -651 -105 -648 -99
rect -660 -108 -648 -105
rect -612 -75 -600 -33
rect -612 -81 -609 -75
rect -603 -81 -600 -75
rect -612 -87 -600 -81
rect -612 -93 -609 -87
rect -603 -93 -600 -87
rect -612 -99 -600 -93
rect -612 -105 -609 -99
rect -603 -105 -600 -99
rect -708 -129 -705 -123
rect -699 -129 -696 -123
rect -708 -132 -696 -129
rect -612 -123 -600 -105
rect -612 -129 -609 -123
rect -603 -129 -600 -123
rect -612 -132 -600 -129
<< via2 >>
rect -705 531 -699 537
rect -657 531 -651 537
rect -705 507 -699 513
rect -705 495 -699 501
rect -705 483 -699 489
rect -609 531 -603 537
rect -657 507 -651 513
rect -657 495 -651 501
rect -657 483 -651 489
rect -657 459 -651 465
rect -681 435 -675 441
rect -705 387 -699 393
rect -609 507 -603 513
rect -609 495 -603 501
rect -609 483 -603 489
rect -633 435 -627 441
rect -681 387 -675 393
rect -657 387 -651 393
rect -633 387 -627 393
rect -609 387 -603 393
rect -681 303 -675 309
rect -705 279 -699 285
rect -705 255 -699 261
rect -705 159 -699 165
rect -705 111 -699 117
rect -705 63 -699 69
rect -705 -33 -699 -27
rect -681 -57 -675 -51
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -633 303 -627 309
rect -609 279 -603 285
rect -609 255 -603 261
rect -609 159 -603 165
rect -609 111 -603 117
rect -609 63 -603 69
rect -609 -33 -603 -27
rect -633 -57 -627 -51
rect -609 -81 -603 -75
rect -609 -93 -603 -87
rect -609 -105 -603 -99
rect -705 -129 -699 -123
rect -609 -129 -603 -123
<< metal3 >>
rect -720 537 -588 540
rect -720 531 -705 537
rect -699 531 -657 537
rect -651 531 -609 537
rect -603 531 -588 537
rect -720 513 -588 531
rect -720 507 -705 513
rect -699 507 -657 513
rect -651 507 -609 513
rect -603 507 -588 513
rect -720 501 -588 507
rect -720 495 -705 501
rect -699 495 -657 501
rect -651 495 -609 501
rect -603 495 -588 501
rect -720 489 -588 495
rect -720 483 -705 489
rect -699 483 -657 489
rect -651 483 -609 489
rect -603 483 -588 489
rect -720 480 -588 483
rect -660 465 -648 468
rect -660 459 -657 465
rect -651 459 -648 465
rect -660 456 -648 459
rect -720 441 -588 444
rect -720 435 -681 441
rect -675 435 -633 441
rect -627 435 -588 441
rect -720 426 -588 435
rect -720 417 -588 420
rect -720 411 -657 417
rect -651 411 -588 417
rect -720 408 -588 411
rect -720 393 -588 402
rect -720 387 -705 393
rect -699 387 -681 393
rect -675 387 -657 393
rect -651 387 -633 393
rect -627 387 -609 393
rect -603 387 -588 393
rect -720 384 -588 387
rect -684 309 -672 312
rect -684 303 -681 309
rect -675 303 -672 309
rect -684 300 -672 303
rect -636 309 -624 312
rect -636 303 -633 309
rect -627 303 -624 309
rect -636 300 -624 303
rect -720 285 -588 288
rect -720 279 -705 285
rect -699 279 -609 285
rect -603 279 -588 285
rect -720 276 -588 279
rect -720 261 -588 264
rect -720 255 -705 261
rect -699 255 -609 261
rect -603 255 -588 261
rect -720 252 -588 255
rect -720 180 -588 240
rect -720 165 -588 168
rect -720 159 -705 165
rect -699 159 -609 165
rect -603 159 -588 165
rect -720 156 -588 159
rect -720 132 -588 144
rect -720 117 -588 120
rect -720 111 -705 117
rect -699 111 -609 117
rect -603 111 -588 117
rect -720 108 -588 111
rect -720 84 -588 96
rect -720 69 -588 72
rect -720 63 -705 69
rect -699 63 -609 69
rect -603 63 -588 69
rect -720 60 -588 63
rect -720 -12 -588 48
rect -720 -27 -588 -24
rect -720 -33 -705 -27
rect -699 -33 -609 -27
rect -603 -33 -588 -27
rect -720 -36 -588 -33
rect -684 -51 -672 -48
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 -51 -624 -48
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
rect -720 -75 -588 -72
rect -720 -81 -705 -75
rect -699 -81 -609 -75
rect -603 -81 -588 -75
rect -720 -87 -588 -81
rect -720 -93 -705 -87
rect -699 -93 -609 -87
rect -603 -93 -588 -87
rect -720 -99 -588 -93
rect -720 -105 -705 -99
rect -699 -105 -609 -99
rect -603 -105 -588 -99
rect -720 -123 -588 -105
rect -720 -129 -705 -123
rect -699 -129 -609 -123
rect -603 -129 -588 -123
rect -720 -132 -588 -129
<< via3 >>
rect -657 459 -651 465
rect -681 435 -675 441
rect -633 435 -627 441
rect -657 411 -651 417
rect -705 387 -699 393
rect -681 387 -675 393
rect -633 387 -627 393
rect -609 387 -603 393
rect -681 303 -675 309
rect -633 303 -627 309
rect -681 -57 -675 -51
rect -633 -57 -627 -51
<< metal4 >>
rect -660 465 -648 468
rect -660 459 -657 465
rect -651 459 -648 465
rect -684 441 -672 444
rect -684 435 -681 441
rect -675 435 -672 441
rect -708 393 -696 396
rect -708 387 -705 393
rect -699 387 -696 393
rect -708 384 -696 387
rect -684 393 -672 435
rect -660 417 -648 459
rect -660 411 -657 417
rect -651 411 -648 417
rect -660 408 -648 411
rect -636 441 -624 444
rect -636 435 -633 441
rect -627 435 -624 441
rect -684 387 -681 393
rect -675 387 -672 393
rect -684 384 -672 387
rect -636 393 -624 435
rect -636 387 -633 393
rect -627 387 -624 393
rect -636 384 -624 387
rect -612 393 -600 396
rect -612 387 -609 393
rect -603 387 -600 393
rect -612 384 -600 387
rect -684 309 -672 312
rect -684 303 -681 309
rect -675 303 -672 309
rect -684 288 -672 303
rect -708 276 -672 288
rect -684 -51 -672 276
rect -684 -57 -681 -51
rect -675 -57 -672 -51
rect -684 -60 -672 -57
rect -636 309 -624 312
rect -636 303 -633 309
rect -627 303 -624 309
rect -636 288 -624 303
rect -636 276 -600 288
rect -636 -51 -624 276
rect -636 -57 -633 -51
rect -627 -57 -624 -51
rect -636 -60 -624 -57
<< labels >>
rlabel metal4 -684 -12 -672 240 0 inl
port 1 nsew
rlabel metal4 -636 -12 -624 240 0 inr
port 2 nsew
rlabel metal2 -660 -12 -648 240 0 out
port 3 nsew
rlabel metal3 -720 480 -588 540 0 vdd
port 4 nsew
rlabel metal3 -720 408 -708 420 0 gp
port 5 nsew
rlabel metal3 -720 276 -708 288 0 bp
port 6 nsew
rlabel metal3 -720 432 -708 444 0 vreg
port 7 nsew
rlabel metal3 -720 180 -588 240 0 op
port 8 nsew
rlabel metal3 -720 132 -588 144 0 im
port 9 nsew
rlabel metal3 -720 84 -588 96 0 ip
port 10 nsew
rlabel metal3 -720 -12 -588 48 0 om
port 11 nsew
rlabel metal3 -720 -132 -588 -72 0 gnd
port 12 nsew
rlabel metal1 -684 -108 -672 -72 0 dl
rlabel metal1 -636 -108 -624 -72 0 dr
rlabel metal1 -708 408 -696 420 0 gnd
rlabel metal1 -708 552 -696 564 0 gnd
<< end >>
