magic
tech gf180mcuC
timestamp 1663277675
<< nwell >>
rect -738 426 -660 546
rect -738 270 -660 402
<< nmos >>
rect -696 -108 -684 -72
<< pmos >>
rect -696 324 -684 354
<< mvpmos >>
rect -696 480 -684 516
<< ndiff >>
rect -708 -75 -696 -72
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
<< pdiff >>
rect -708 345 -696 354
rect -708 339 -705 345
rect -699 339 -696 345
rect -708 333 -696 339
rect -708 327 -705 333
rect -699 327 -696 333
rect -708 324 -696 327
rect -684 345 -672 354
rect -684 339 -681 345
rect -675 339 -672 345
rect -684 333 -672 339
rect -684 327 -681 333
rect -675 327 -672 333
rect -684 324 -672 327
<< mvpdiff >>
rect -708 513 -696 516
rect -708 507 -705 513
rect -699 507 -696 513
rect -708 501 -696 507
rect -708 495 -705 501
rect -699 495 -696 501
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 480 -696 483
rect -684 513 -672 516
rect -684 507 -681 513
rect -675 507 -672 513
rect -684 501 -672 507
rect -684 495 -681 501
rect -675 495 -672 501
rect -684 489 -672 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
<< ndiffc >>
rect -705 -81 -699 -75
rect -705 -93 -699 -87
rect -705 -105 -699 -99
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
<< pdiffc >>
rect -705 339 -699 345
rect -705 327 -699 333
rect -681 339 -675 345
rect -681 327 -675 333
<< mvpdiffc >>
rect -705 507 -699 513
rect -705 495 -699 501
rect -705 483 -699 489
rect -681 507 -675 513
rect -681 495 -675 501
rect -681 483 -675 489
<< psubdiff >>
rect -756 561 -660 564
rect -756 555 -753 561
rect -747 555 -741 561
rect -735 555 -729 561
rect -723 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -660 561
rect -756 552 -660 555
rect -756 549 -744 552
rect -756 543 -753 549
rect -747 543 -744 549
rect -756 537 -744 543
rect -756 531 -753 537
rect -747 531 -744 537
rect -756 525 -744 531
rect -756 519 -753 525
rect -747 519 -744 525
rect -756 513 -744 519
rect -756 507 -753 513
rect -747 507 -744 513
rect -756 501 -744 507
rect -756 495 -753 501
rect -747 495 -744 501
rect -756 489 -744 495
rect -756 483 -753 489
rect -747 483 -744 489
rect -756 477 -744 483
rect -756 471 -753 477
rect -747 471 -744 477
rect -756 465 -744 471
rect -756 459 -753 465
rect -747 459 -744 465
rect -756 453 -744 459
rect -756 447 -753 453
rect -747 447 -744 453
rect -756 441 -744 447
rect -756 435 -753 441
rect -747 435 -744 441
rect -756 429 -744 435
rect -756 423 -753 429
rect -747 423 -744 429
rect -756 420 -744 423
rect -756 417 -660 420
rect -756 411 -753 417
rect -747 411 -741 417
rect -735 411 -729 417
rect -723 411 -717 417
rect -711 411 -705 417
rect -699 411 -693 417
rect -687 411 -681 417
rect -675 411 -669 417
rect -663 411 -660 417
rect -756 408 -660 411
rect -756 405 -744 408
rect -756 399 -753 405
rect -747 399 -744 405
rect -756 393 -744 399
rect -756 387 -753 393
rect -747 387 -744 393
rect -756 381 -744 387
rect -756 375 -753 381
rect -747 375 -744 381
rect -756 369 -744 375
rect -756 363 -753 369
rect -747 363 -744 369
rect -756 357 -744 363
rect -756 351 -753 357
rect -747 351 -744 357
rect -756 345 -744 351
rect -756 339 -753 345
rect -747 339 -744 345
rect -756 333 -744 339
rect -756 327 -753 333
rect -747 327 -744 333
rect -756 321 -744 327
rect -756 315 -753 321
rect -747 315 -744 321
rect -756 309 -744 315
rect -756 303 -753 309
rect -747 303 -744 309
rect -756 297 -744 303
rect -756 291 -753 297
rect -747 291 -744 297
rect -756 285 -744 291
rect -756 279 -753 285
rect -747 279 -744 285
rect -756 273 -744 279
rect -756 267 -753 273
rect -747 267 -744 273
rect -756 264 -744 267
rect -756 261 -660 264
rect -756 255 -753 261
rect -747 255 -741 261
rect -735 255 -729 261
rect -723 255 -717 261
rect -711 255 -705 261
rect -699 255 -693 261
rect -687 255 -681 261
rect -675 255 -669 261
rect -663 255 -660 261
rect -756 252 -660 255
rect -756 249 -744 252
rect -756 243 -753 249
rect -747 243 -744 249
rect -756 237 -744 243
rect -756 231 -753 237
rect -747 231 -744 237
rect -756 225 -744 231
rect -756 219 -753 225
rect -747 219 -744 225
rect -756 213 -744 219
rect -756 207 -753 213
rect -747 207 -744 213
rect -756 201 -744 207
rect -756 195 -753 201
rect -747 195 -744 201
rect -756 189 -744 195
rect -756 183 -753 189
rect -747 183 -744 189
rect -756 177 -744 183
rect -756 171 -753 177
rect -747 171 -744 177
rect -756 168 -744 171
rect -756 165 -660 168
rect -756 159 -753 165
rect -747 159 -741 165
rect -735 159 -729 165
rect -723 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -660 165
rect -756 156 -660 159
rect -756 153 -744 156
rect -756 147 -753 153
rect -747 147 -744 153
rect -756 141 -744 147
rect -756 135 -753 141
rect -747 135 -744 141
rect -756 129 -744 135
rect -756 123 -753 129
rect -747 123 -744 129
rect -756 120 -744 123
rect -756 117 -660 120
rect -756 111 -753 117
rect -747 111 -741 117
rect -735 111 -729 117
rect -723 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -660 117
rect -756 108 -660 111
rect -756 105 -744 108
rect -756 99 -753 105
rect -747 99 -744 105
rect -756 93 -744 99
rect -756 87 -753 93
rect -747 87 -744 93
rect -756 81 -744 87
rect -756 75 -753 81
rect -747 75 -744 81
rect -756 72 -744 75
rect -756 69 -660 72
rect -756 63 -753 69
rect -747 63 -741 69
rect -735 63 -729 69
rect -723 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -660 69
rect -756 60 -660 63
rect -756 57 -744 60
rect -756 51 -753 57
rect -747 51 -744 57
rect -756 45 -744 51
rect -756 39 -753 45
rect -747 39 -744 45
rect -756 33 -744 39
rect -756 27 -753 33
rect -747 27 -744 33
rect -756 21 -744 27
rect -756 15 -753 21
rect -747 15 -744 21
rect -756 9 -744 15
rect -756 3 -753 9
rect -747 3 -744 9
rect -756 -3 -744 3
rect -756 -9 -753 -3
rect -747 -9 -744 -3
rect -756 -15 -744 -9
rect -756 -21 -753 -15
rect -747 -21 -744 -15
rect -756 -24 -744 -21
rect -756 -27 -660 -24
rect -756 -33 -753 -27
rect -747 -33 -741 -27
rect -735 -33 -729 -27
rect -723 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -39 -744 -36
rect -756 -45 -753 -39
rect -747 -45 -744 -39
rect -756 -51 -744 -45
rect -756 -57 -753 -51
rect -747 -57 -744 -51
rect -756 -63 -744 -57
rect -756 -69 -753 -63
rect -747 -69 -744 -63
rect -756 -75 -744 -69
rect -756 -81 -753 -75
rect -747 -81 -744 -75
rect -756 -87 -744 -81
rect -756 -93 -753 -87
rect -747 -93 -744 -87
rect -756 -99 -744 -93
rect -756 -105 -753 -99
rect -747 -105 -744 -99
rect -756 -111 -744 -105
rect -756 -117 -753 -111
rect -747 -117 -744 -111
rect -756 -120 -744 -117
rect -756 -123 -660 -120
rect -756 -129 -753 -123
rect -747 -129 -741 -123
rect -735 -129 -729 -123
rect -723 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -660 -123
rect -756 -132 -660 -129
<< nsubdiff >>
rect -732 393 -672 396
rect -732 387 -729 393
rect -723 387 -717 393
rect -711 387 -705 393
rect -699 387 -693 393
rect -687 387 -681 393
rect -675 387 -672 393
rect -732 384 -672 387
rect -732 381 -720 384
rect -732 375 -729 381
rect -723 375 -720 381
rect -732 369 -720 375
rect -732 363 -729 369
rect -723 363 -720 369
rect -732 357 -720 363
rect -732 351 -729 357
rect -723 351 -720 357
rect -732 345 -720 351
rect -732 339 -729 345
rect -723 339 -720 345
rect -732 333 -720 339
rect -732 327 -729 333
rect -723 327 -720 333
rect -732 321 -720 327
rect -732 315 -729 321
rect -723 315 -720 321
rect -732 309 -720 315
rect -732 303 -729 309
rect -723 303 -720 309
rect -732 297 -720 303
rect -732 291 -729 297
rect -723 291 -720 297
rect -732 288 -720 291
rect -732 285 -672 288
rect -732 279 -729 285
rect -723 279 -717 285
rect -711 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -672 285
rect -732 276 -672 279
<< mvnsubdiff >>
rect -732 537 -672 540
rect -732 531 -729 537
rect -723 531 -717 537
rect -711 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -672 537
rect -732 528 -672 531
rect -732 525 -720 528
rect -732 519 -729 525
rect -723 519 -720 525
rect -732 513 -720 519
rect -732 507 -729 513
rect -723 507 -720 513
rect -732 501 -720 507
rect -732 495 -729 501
rect -723 495 -720 501
rect -732 489 -720 495
rect -732 483 -729 489
rect -723 483 -720 489
rect -732 477 -720 483
rect -732 471 -729 477
rect -723 471 -720 477
rect -732 465 -720 471
rect -732 459 -729 465
rect -723 459 -720 465
rect -732 453 -720 459
rect -732 447 -729 453
rect -723 447 -720 453
rect -732 444 -720 447
rect -732 441 -672 444
rect -732 435 -729 441
rect -723 435 -717 441
rect -711 435 -705 441
rect -699 435 -693 441
rect -687 435 -681 441
rect -675 435 -672 441
rect -732 432 -672 435
<< psubdiffcont >>
rect -753 555 -747 561
rect -741 555 -735 561
rect -729 555 -723 561
rect -717 555 -711 561
rect -705 555 -699 561
rect -693 555 -687 561
rect -681 555 -675 561
rect -669 555 -663 561
rect -753 543 -747 549
rect -753 531 -747 537
rect -753 519 -747 525
rect -753 507 -747 513
rect -753 495 -747 501
rect -753 483 -747 489
rect -753 471 -747 477
rect -753 459 -747 465
rect -753 447 -747 453
rect -753 435 -747 441
rect -753 423 -747 429
rect -753 411 -747 417
rect -741 411 -735 417
rect -729 411 -723 417
rect -717 411 -711 417
rect -705 411 -699 417
rect -693 411 -687 417
rect -681 411 -675 417
rect -669 411 -663 417
rect -753 399 -747 405
rect -753 387 -747 393
rect -753 375 -747 381
rect -753 363 -747 369
rect -753 351 -747 357
rect -753 339 -747 345
rect -753 327 -747 333
rect -753 315 -747 321
rect -753 303 -747 309
rect -753 291 -747 297
rect -753 279 -747 285
rect -753 267 -747 273
rect -753 255 -747 261
rect -741 255 -735 261
rect -729 255 -723 261
rect -717 255 -711 261
rect -705 255 -699 261
rect -693 255 -687 261
rect -681 255 -675 261
rect -669 255 -663 261
rect -753 243 -747 249
rect -753 231 -747 237
rect -753 219 -747 225
rect -753 207 -747 213
rect -753 195 -747 201
rect -753 183 -747 189
rect -753 171 -747 177
rect -753 159 -747 165
rect -741 159 -735 165
rect -729 159 -723 165
rect -717 159 -711 165
rect -705 159 -699 165
rect -693 159 -687 165
rect -681 159 -675 165
rect -669 159 -663 165
rect -753 147 -747 153
rect -753 135 -747 141
rect -753 123 -747 129
rect -753 111 -747 117
rect -741 111 -735 117
rect -729 111 -723 117
rect -717 111 -711 117
rect -705 111 -699 117
rect -693 111 -687 117
rect -681 111 -675 117
rect -669 111 -663 117
rect -753 99 -747 105
rect -753 87 -747 93
rect -753 75 -747 81
rect -753 63 -747 69
rect -741 63 -735 69
rect -729 63 -723 69
rect -717 63 -711 69
rect -705 63 -699 69
rect -693 63 -687 69
rect -681 63 -675 69
rect -669 63 -663 69
rect -753 51 -747 57
rect -753 39 -747 45
rect -753 27 -747 33
rect -753 15 -747 21
rect -753 3 -747 9
rect -753 -9 -747 -3
rect -753 -21 -747 -15
rect -753 -33 -747 -27
rect -741 -33 -735 -27
rect -729 -33 -723 -27
rect -717 -33 -711 -27
rect -705 -33 -699 -27
rect -693 -33 -687 -27
rect -681 -33 -675 -27
rect -669 -33 -663 -27
rect -753 -45 -747 -39
rect -753 -57 -747 -51
rect -753 -69 -747 -63
rect -753 -81 -747 -75
rect -753 -93 -747 -87
rect -753 -105 -747 -99
rect -753 -117 -747 -111
rect -753 -129 -747 -123
rect -741 -129 -735 -123
rect -729 -129 -723 -123
rect -717 -129 -711 -123
rect -705 -129 -699 -123
rect -693 -129 -687 -123
rect -681 -129 -675 -123
rect -669 -129 -663 -123
<< nsubdiffcont >>
rect -729 387 -723 393
rect -717 387 -711 393
rect -705 387 -699 393
rect -693 387 -687 393
rect -681 387 -675 393
rect -729 375 -723 381
rect -729 363 -723 369
rect -729 351 -723 357
rect -729 339 -723 345
rect -729 327 -723 333
rect -729 315 -723 321
rect -729 303 -723 309
rect -729 291 -723 297
rect -729 279 -723 285
rect -717 279 -711 285
rect -705 279 -699 285
rect -693 279 -687 285
rect -681 279 -675 285
<< mvnsubdiffcont >>
rect -729 531 -723 537
rect -717 531 -711 537
rect -705 531 -699 537
rect -693 531 -687 537
rect -681 531 -675 537
rect -729 519 -723 525
rect -729 507 -723 513
rect -729 495 -723 501
rect -729 483 -723 489
rect -729 471 -723 477
rect -729 459 -723 465
rect -729 447 -723 453
rect -729 435 -723 441
rect -717 435 -711 441
rect -705 435 -699 441
rect -693 435 -687 441
rect -681 435 -675 441
<< polysilicon >>
rect -696 516 -684 522
rect -696 465 -684 480
rect -696 459 -693 465
rect -687 459 -684 465
rect -696 456 -684 459
rect -696 354 -684 360
rect -696 309 -684 324
rect -696 303 -693 309
rect -687 303 -684 309
rect -696 300 -684 303
rect -696 -51 -684 -48
rect -696 -57 -693 -51
rect -687 -57 -684 -51
rect -696 -72 -684 -57
rect -696 -114 -684 -108
<< polycontact >>
rect -693 459 -687 465
rect -693 303 -687 309
rect -693 -57 -687 -51
<< metal1 >>
rect -756 561 -660 564
rect -756 555 -753 561
rect -747 555 -741 561
rect -735 555 -729 561
rect -723 555 -717 561
rect -711 555 -705 561
rect -699 555 -693 561
rect -687 555 -681 561
rect -675 555 -669 561
rect -663 555 -660 561
rect -756 552 -660 555
rect -756 549 -744 552
rect -756 543 -753 549
rect -747 543 -744 549
rect -756 537 -744 543
rect -756 531 -753 537
rect -747 531 -744 537
rect -756 525 -744 531
rect -756 519 -753 525
rect -747 519 -744 525
rect -756 513 -744 519
rect -756 507 -753 513
rect -747 507 -744 513
rect -756 501 -744 507
rect -756 495 -753 501
rect -747 495 -744 501
rect -756 489 -744 495
rect -756 483 -753 489
rect -747 483 -744 489
rect -756 477 -744 483
rect -756 471 -753 477
rect -747 471 -744 477
rect -756 465 -744 471
rect -756 459 -753 465
rect -747 459 -744 465
rect -756 453 -744 459
rect -756 447 -753 453
rect -747 447 -744 453
rect -756 441 -744 447
rect -756 435 -753 441
rect -747 435 -744 441
rect -756 429 -744 435
rect -732 537 -660 540
rect -732 531 -729 537
rect -723 531 -717 537
rect -711 531 -705 537
rect -699 531 -693 537
rect -687 531 -681 537
rect -675 531 -660 537
rect -732 528 -660 531
rect -732 525 -720 528
rect -732 519 -729 525
rect -723 519 -720 525
rect -732 513 -720 519
rect -732 507 -729 513
rect -723 507 -720 513
rect -732 501 -720 507
rect -732 495 -729 501
rect -723 495 -720 501
rect -732 489 -720 495
rect -732 483 -729 489
rect -723 483 -720 489
rect -732 477 -720 483
rect -732 471 -729 477
rect -723 471 -720 477
rect -732 465 -720 471
rect -732 459 -729 465
rect -723 459 -720 465
rect -732 453 -720 459
rect -708 513 -696 516
rect -708 507 -705 513
rect -699 507 -696 513
rect -708 501 -696 507
rect -708 495 -705 501
rect -699 495 -696 501
rect -708 489 -696 495
rect -708 483 -705 489
rect -699 483 -696 489
rect -708 468 -696 483
rect -684 513 -672 516
rect -684 507 -681 513
rect -675 507 -672 513
rect -684 501 -672 507
rect -684 495 -681 501
rect -675 495 -672 501
rect -684 489 -672 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -708 465 -684 468
rect -708 459 -693 465
rect -687 459 -684 465
rect -708 456 -684 459
rect -732 447 -729 453
rect -723 447 -720 453
rect -732 444 -720 447
rect -732 441 -660 444
rect -732 435 -729 441
rect -723 435 -717 441
rect -711 435 -705 441
rect -699 435 -693 441
rect -687 435 -681 441
rect -675 435 -660 441
rect -732 432 -660 435
rect -756 423 -753 429
rect -747 423 -744 429
rect -756 420 -744 423
rect -756 417 -660 420
rect -756 411 -753 417
rect -747 411 -741 417
rect -735 411 -729 417
rect -723 411 -717 417
rect -711 411 -705 417
rect -699 411 -693 417
rect -687 411 -681 417
rect -675 411 -669 417
rect -663 411 -660 417
rect -756 408 -660 411
rect -756 405 -744 408
rect -756 399 -753 405
rect -747 399 -744 405
rect -756 393 -744 399
rect -756 387 -753 393
rect -747 387 -744 393
rect -756 381 -744 387
rect -756 375 -753 381
rect -747 375 -744 381
rect -756 369 -744 375
rect -756 363 -753 369
rect -747 363 -744 369
rect -756 357 -744 363
rect -756 351 -753 357
rect -747 351 -744 357
rect -756 345 -744 351
rect -756 339 -753 345
rect -747 339 -744 345
rect -756 333 -744 339
rect -756 327 -753 333
rect -747 327 -744 333
rect -756 321 -744 327
rect -756 315 -753 321
rect -747 315 -744 321
rect -756 309 -744 315
rect -756 303 -753 309
rect -747 303 -744 309
rect -756 297 -744 303
rect -756 291 -753 297
rect -747 291 -744 297
rect -756 285 -744 291
rect -756 279 -753 285
rect -747 279 -744 285
rect -756 273 -744 279
rect -732 393 -672 396
rect -732 387 -729 393
rect -723 387 -717 393
rect -711 387 -705 393
rect -699 387 -693 393
rect -687 387 -681 393
rect -675 387 -672 393
rect -732 384 -672 387
rect -732 381 -720 384
rect -732 375 -729 381
rect -723 375 -720 381
rect -732 369 -720 375
rect -732 363 -729 369
rect -723 363 -720 369
rect -732 357 -720 363
rect -732 351 -729 357
rect -723 351 -720 357
rect -732 345 -720 351
rect -732 339 -729 345
rect -723 339 -720 345
rect -732 333 -720 339
rect -732 327 -729 333
rect -723 327 -720 333
rect -732 321 -720 327
rect -732 315 -729 321
rect -723 315 -720 321
rect -732 309 -720 315
rect -732 303 -729 309
rect -723 303 -720 309
rect -732 297 -720 303
rect -708 345 -696 354
rect -708 339 -705 345
rect -699 339 -696 345
rect -708 333 -696 339
rect -708 327 -705 333
rect -699 327 -696 333
rect -708 312 -696 327
rect -684 345 -672 354
rect -684 339 -681 345
rect -675 339 -672 345
rect -684 333 -672 339
rect -684 327 -681 333
rect -675 327 -672 333
rect -684 324 -672 327
rect -708 309 -684 312
rect -708 303 -693 309
rect -687 303 -684 309
rect -708 300 -684 303
rect -732 291 -729 297
rect -723 291 -720 297
rect -732 288 -720 291
rect -732 285 -660 288
rect -732 279 -729 285
rect -723 279 -717 285
rect -711 279 -705 285
rect -699 279 -693 285
rect -687 279 -681 285
rect -675 279 -660 285
rect -732 276 -660 279
rect -756 267 -753 273
rect -747 267 -744 273
rect -756 264 -744 267
rect -756 261 -660 264
rect -756 255 -753 261
rect -747 255 -741 261
rect -735 255 -729 261
rect -723 255 -717 261
rect -711 255 -705 261
rect -699 255 -693 261
rect -687 255 -681 261
rect -675 255 -669 261
rect -663 255 -660 261
rect -756 252 -660 255
rect -756 249 -744 252
rect -756 243 -753 249
rect -747 243 -744 249
rect -756 237 -744 243
rect -756 231 -753 237
rect -747 231 -744 237
rect -756 225 -744 231
rect -756 219 -753 225
rect -747 219 -744 225
rect -756 213 -744 219
rect -756 207 -753 213
rect -747 207 -744 213
rect -756 201 -744 207
rect -756 195 -753 201
rect -747 195 -744 201
rect -756 189 -744 195
rect -756 183 -753 189
rect -747 183 -744 189
rect -756 177 -744 183
rect -756 171 -753 177
rect -747 171 -744 177
rect -756 168 -744 171
rect -756 165 -660 168
rect -756 159 -753 165
rect -747 159 -741 165
rect -735 159 -729 165
rect -723 159 -717 165
rect -711 159 -705 165
rect -699 159 -693 165
rect -687 159 -681 165
rect -675 159 -669 165
rect -663 159 -660 165
rect -756 156 -660 159
rect -756 153 -744 156
rect -756 147 -753 153
rect -747 147 -744 153
rect -756 141 -744 147
rect -756 135 -753 141
rect -747 135 -744 141
rect -756 129 -744 135
rect -756 123 -753 129
rect -747 123 -744 129
rect -756 120 -744 123
rect -756 117 -660 120
rect -756 111 -753 117
rect -747 111 -741 117
rect -735 111 -729 117
rect -723 111 -717 117
rect -711 111 -705 117
rect -699 111 -693 117
rect -687 111 -681 117
rect -675 111 -669 117
rect -663 111 -660 117
rect -756 108 -660 111
rect -756 105 -744 108
rect -756 99 -753 105
rect -747 99 -744 105
rect -756 93 -744 99
rect -756 87 -753 93
rect -747 87 -744 93
rect -756 81 -744 87
rect -756 75 -753 81
rect -747 75 -744 81
rect -756 72 -744 75
rect -756 69 -660 72
rect -756 63 -753 69
rect -747 63 -741 69
rect -735 63 -729 69
rect -723 63 -717 69
rect -711 63 -705 69
rect -699 63 -693 69
rect -687 63 -681 69
rect -675 63 -669 69
rect -663 63 -660 69
rect -756 60 -660 63
rect -756 57 -744 60
rect -756 51 -753 57
rect -747 51 -744 57
rect -756 45 -744 51
rect -756 39 -753 45
rect -747 39 -744 45
rect -756 33 -744 39
rect -756 27 -753 33
rect -747 27 -744 33
rect -756 21 -744 27
rect -756 15 -753 21
rect -747 15 -744 21
rect -756 9 -744 15
rect -756 3 -753 9
rect -747 3 -744 9
rect -756 -3 -744 3
rect -756 -9 -753 -3
rect -747 -9 -744 -3
rect -756 -15 -744 -9
rect -756 -21 -753 -15
rect -747 -21 -744 -15
rect -756 -24 -744 -21
rect -756 -27 -660 -24
rect -756 -33 -753 -27
rect -747 -33 -741 -27
rect -735 -33 -729 -27
rect -723 -33 -717 -27
rect -711 -33 -705 -27
rect -699 -33 -693 -27
rect -687 -33 -681 -27
rect -675 -33 -669 -27
rect -663 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -39 -744 -36
rect -756 -45 -753 -39
rect -747 -45 -744 -39
rect -756 -51 -744 -45
rect -756 -57 -753 -51
rect -747 -57 -744 -51
rect -756 -63 -744 -57
rect -756 -69 -753 -63
rect -747 -69 -744 -63
rect -756 -75 -744 -69
rect -756 -81 -753 -75
rect -747 -81 -744 -75
rect -756 -87 -744 -81
rect -756 -93 -753 -87
rect -747 -93 -744 -87
rect -756 -99 -744 -93
rect -756 -105 -753 -99
rect -747 -105 -744 -99
rect -756 -111 -744 -105
rect -708 -51 -684 -48
rect -708 -57 -693 -51
rect -687 -57 -684 -51
rect -708 -60 -684 -57
rect -708 -75 -696 -60
rect -708 -81 -705 -75
rect -699 -81 -696 -75
rect -708 -87 -696 -81
rect -708 -93 -705 -87
rect -699 -93 -696 -87
rect -708 -99 -696 -93
rect -708 -105 -705 -99
rect -699 -105 -696 -99
rect -708 -108 -696 -105
rect -684 -75 -672 -72
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -108 -672 -105
rect -756 -117 -753 -111
rect -747 -117 -744 -111
rect -756 -120 -744 -117
rect -756 -123 -660 -120
rect -756 -129 -753 -123
rect -747 -129 -741 -123
rect -735 -129 -729 -123
rect -723 -129 -717 -123
rect -711 -129 -705 -123
rect -699 -129 -693 -123
rect -687 -129 -681 -123
rect -675 -129 -669 -123
rect -663 -129 -660 -123
rect -756 -132 -660 -129
<< via1 >>
rect -681 531 -675 537
rect -681 507 -675 513
rect -681 495 -675 501
rect -681 483 -675 489
rect -681 339 -675 345
rect -681 327 -675 333
rect -729 279 -723 285
rect -681 255 -675 261
rect -681 159 -675 165
rect -681 111 -675 117
rect -681 63 -675 69
rect -681 -33 -675 -27
rect -681 -81 -675 -75
rect -681 -93 -675 -87
rect -681 -105 -675 -99
rect -681 -129 -675 -123
<< metal2 >>
rect -684 537 -672 540
rect -684 531 -681 537
rect -675 531 -672 537
rect -684 513 -672 531
rect -684 507 -681 513
rect -675 507 -672 513
rect -684 501 -672 507
rect -684 495 -681 501
rect -675 495 -672 501
rect -684 489 -672 495
rect -684 483 -681 489
rect -675 483 -672 489
rect -684 480 -672 483
rect -708 441 -696 444
rect -708 435 -705 441
rect -699 435 -696 441
rect -708 393 -696 435
rect -708 387 -705 393
rect -699 387 -696 393
rect -708 384 -696 387
rect -684 393 -672 396
rect -684 387 -681 393
rect -675 387 -672 393
rect -684 345 -672 387
rect -684 339 -681 345
rect -675 339 -672 345
rect -684 333 -672 339
rect -684 327 -681 333
rect -675 327 -672 333
rect -684 324 -672 327
rect -732 285 -720 288
rect -732 279 -729 285
rect -723 279 -720 285
rect -732 276 -720 279
rect -684 261 -672 264
rect -684 255 -681 261
rect -675 255 -672 261
rect -684 165 -672 255
rect -684 159 -681 165
rect -675 159 -672 165
rect -684 117 -672 159
rect -684 111 -681 117
rect -675 111 -672 117
rect -684 69 -672 111
rect -684 63 -681 69
rect -675 63 -672 69
rect -684 -27 -672 63
rect -684 -33 -681 -27
rect -675 -33 -672 -27
rect -684 -75 -672 -33
rect -684 -81 -681 -75
rect -675 -81 -672 -75
rect -684 -87 -672 -81
rect -684 -93 -681 -87
rect -675 -93 -672 -87
rect -684 -99 -672 -93
rect -684 -105 -681 -99
rect -675 -105 -672 -99
rect -684 -123 -672 -105
rect -684 -129 -681 -123
rect -675 -129 -672 -123
rect -684 -132 -672 -129
<< via2 >>
rect -681 531 -675 537
rect -681 507 -675 513
rect -681 495 -675 501
rect -681 483 -675 489
rect -705 435 -699 441
rect -705 387 -699 393
rect -681 387 -675 393
rect -729 279 -723 285
rect -681 255 -675 261
rect -681 159 -675 165
rect -681 111 -675 117
rect -681 63 -675 69
rect -681 -33 -675 -27
rect -681 -129 -675 -123
<< metal3 >>
rect -756 537 -660 540
rect -756 531 -681 537
rect -675 531 -660 537
rect -756 513 -660 531
rect -756 507 -681 513
rect -675 507 -660 513
rect -756 501 -660 507
rect -756 495 -681 501
rect -675 495 -660 501
rect -756 489 -660 495
rect -756 483 -681 489
rect -675 483 -660 489
rect -756 480 -660 483
rect -756 441 -660 444
rect -756 435 -705 441
rect -699 435 -660 441
rect -756 426 -660 435
rect -756 408 -660 420
rect -756 393 -660 402
rect -756 387 -705 393
rect -699 387 -681 393
rect -675 387 -660 393
rect -756 384 -660 387
rect -756 285 -660 288
rect -756 279 -729 285
rect -723 279 -660 285
rect -756 276 -660 279
rect -756 261 -660 264
rect -756 255 -681 261
rect -675 255 -660 261
rect -756 252 -660 255
rect -756 180 -660 240
rect -756 165 -660 168
rect -756 159 -681 165
rect -675 159 -660 165
rect -756 156 -660 159
rect -756 132 -660 144
rect -756 117 -660 120
rect -756 111 -681 117
rect -675 111 -660 117
rect -756 108 -660 111
rect -756 84 -660 96
rect -756 69 -660 72
rect -756 63 -681 69
rect -675 63 -660 69
rect -756 60 -660 63
rect -756 -12 -660 48
rect -756 -27 -660 -24
rect -756 -33 -681 -27
rect -675 -33 -660 -27
rect -756 -36 -660 -33
rect -756 -123 -660 -72
rect -756 -129 -681 -123
rect -675 -129 -660 -123
rect -756 -132 -660 -129
<< labels >>
rlabel metal3 -756 480 -660 540 0 vdd
port 1 nsew
rlabel metal3 -756 408 -660 420 0 gp
port 2 nsew
rlabel metal3 -756 276 -660 288 0 bp
port 3 nsew
rlabel metal3 -756 432 -660 444 0 vreg
port 4 nsew
rlabel metal3 -756 180 -660 240 0 op
port 5 nsew
rlabel metal3 -756 132 -660 144 0 im
port 6 nsew
rlabel metal3 -756 84 -660 96 0 ip
port 7 nsew
rlabel metal3 -756 -12 -660 48 0 om
port 8 nsew
rlabel metal3 -756 -132 -660 -72 0 gnd
port 9 nsew
rlabel metal1 -708 456 -696 468 1 hih
rlabel metal1 -708 300 -696 312 0 hi
rlabel metal1 -708 -60 -696 -48 0 lo
<< end >>
