magic
tech gf180mcuC
timestamp 1665299032
<< via2 >>
rect -768 324 -756 348
rect -648 324 -636 348
rect 792 324 804 348
rect 912 324 924 348
rect 1272 324 1284 348
rect 1392 324 1404 348
rect 2832 324 2844 348
rect 2952 324 2964 348
rect -288 300 -276 312
rect 432 300 444 312
rect 1752 300 1764 312
rect 2472 300 2484 312
rect -768 264 -756 288
rect -648 264 -636 288
rect 792 264 804 288
rect 912 264 924 288
rect 1272 264 1284 288
rect 1392 264 1404 288
rect 2832 264 2844 288
rect 2952 264 2964 288
rect -168 168 -156 180
rect 312 168 324 180
rect 1872 168 1884 180
rect 2352 168 2364 180
rect -48 120 -36 132
rect 72 120 84 132
rect 192 120 204 132
rect 1992 120 2004 132
rect 2112 120 2124 132
rect 2232 120 2244 132
rect -888 12 -876 36
rect -528 12 -516 36
rect 672 12 684 36
rect 1032 12 1044 36
rect 1152 12 1164 36
rect 1512 12 1524 36
rect 2712 12 2724 36
rect 3072 12 3084 36
rect -408 -12 -396 0
rect 552 -12 564 0
rect 1632 -12 1644 0
rect 2592 -12 2604 0
rect -888 -48 -876 -24
rect -528 -48 -516 -24
rect 672 -48 684 -24
rect 1032 -48 1044 -24
rect 1152 -48 1164 -24
rect 1512 -48 1524 -24
rect 2712 -48 2724 -24
rect 3072 -48 3084 -24
<< mimcap >>
rect -1008 876 2976 888
rect -1008 864 -996 876
rect -984 864 -948 876
rect -936 864 -924 876
rect -912 864 -876 876
rect -864 864 -852 876
rect -840 864 -804 876
rect -792 864 -780 876
rect -768 864 -732 876
rect -720 864 -708 876
rect -696 864 -660 876
rect -648 864 -636 876
rect -624 864 -588 876
rect -576 864 -564 876
rect -552 864 -516 876
rect -504 864 -492 876
rect -480 864 -444 876
rect -432 864 -420 876
rect -408 864 -372 876
rect -360 864 -348 876
rect -336 864 -300 876
rect -288 864 -276 876
rect -264 864 -228 876
rect -216 864 -204 876
rect -192 864 -156 876
rect -144 864 -132 876
rect -120 864 -84 876
rect -72 864 -60 876
rect -48 864 -12 876
rect 0 864 12 876
rect 24 864 60 876
rect 72 864 84 876
rect 96 864 132 876
rect 144 864 156 876
rect 168 864 204 876
rect 216 864 228 876
rect 240 864 276 876
rect 288 864 300 876
rect 312 864 348 876
rect 360 864 372 876
rect 384 864 420 876
rect 432 864 444 876
rect 456 864 492 876
rect 504 864 516 876
rect 528 864 564 876
rect 576 864 588 876
rect 600 864 636 876
rect 648 864 660 876
rect 672 864 708 876
rect 720 864 732 876
rect 744 864 780 876
rect 792 864 804 876
rect 816 864 852 876
rect 864 864 876 876
rect 888 864 924 876
rect 936 864 948 876
rect 960 864 996 876
rect 1008 864 1020 876
rect 1032 864 1068 876
rect 1080 864 1092 876
rect 1104 864 1140 876
rect 1152 864 1164 876
rect 1176 864 1212 876
rect 1224 864 1236 876
rect 1248 864 1284 876
rect 1296 864 1308 876
rect 1320 864 1356 876
rect 1368 864 1380 876
rect 1392 864 1428 876
rect 1440 864 1452 876
rect 1464 864 1500 876
rect 1512 864 1524 876
rect 1536 864 1572 876
rect 1584 864 1596 876
rect 1608 864 1644 876
rect 1656 864 1668 876
rect 1680 864 1716 876
rect 1728 864 1740 876
rect 1752 864 1788 876
rect 1800 864 1812 876
rect 1824 864 1860 876
rect 1872 864 1884 876
rect 1896 864 1932 876
rect 1944 864 1956 876
rect 1968 864 2004 876
rect 2016 864 2028 876
rect 2040 864 2076 876
rect 2088 864 2100 876
rect 2112 864 2148 876
rect 2160 864 2172 876
rect 2184 864 2220 876
rect 2232 864 2244 876
rect 2256 864 2292 876
rect 2304 864 2316 876
rect 2328 864 2364 876
rect 2376 864 2388 876
rect 2400 864 2436 876
rect 2448 864 2460 876
rect 2472 864 2484 876
rect 2496 864 2532 876
rect 2544 864 2556 876
rect 2568 864 2604 876
rect 2616 864 2628 876
rect 2640 864 2676 876
rect 2688 864 2700 876
rect 2712 864 2724 876
rect 2736 864 2772 876
rect 2784 864 2796 876
rect 2808 864 2844 876
rect 2856 864 2868 876
rect 2880 864 2916 876
rect 2928 864 2940 876
rect 2952 864 2976 876
rect -1008 840 2976 864
rect -1008 828 -996 840
rect -984 828 -972 840
rect -960 828 -948 840
rect -936 828 -924 840
rect -912 828 -900 840
rect -888 828 -876 840
rect -864 828 -852 840
rect -840 828 -828 840
rect -816 828 -804 840
rect -792 828 -780 840
rect -768 828 -756 840
rect -744 828 -732 840
rect -720 828 -708 840
rect -696 828 -684 840
rect -672 828 -660 840
rect -648 828 -636 840
rect -624 828 -612 840
rect -600 828 -588 840
rect -576 828 -564 840
rect -552 828 -540 840
rect -528 828 -516 840
rect -504 828 -492 840
rect -480 828 -468 840
rect -456 828 -444 840
rect -432 828 -420 840
rect -408 828 -396 840
rect -384 828 -372 840
rect -360 828 -348 840
rect -336 828 -324 840
rect -312 828 -300 840
rect -288 828 -276 840
rect -264 828 -252 840
rect -240 828 -228 840
rect -216 828 -204 840
rect -192 828 -180 840
rect -168 828 -156 840
rect -144 828 -132 840
rect -120 828 -108 840
rect -96 828 -84 840
rect -72 828 -60 840
rect -48 828 -36 840
rect -24 828 -12 840
rect 0 828 12 840
rect 24 828 36 840
rect 48 828 60 840
rect 72 828 84 840
rect 96 828 108 840
rect 120 828 132 840
rect 144 828 156 840
rect 168 828 180 840
rect 192 828 204 840
rect 216 828 228 840
rect 240 828 252 840
rect 264 828 276 840
rect 288 828 300 840
rect 312 828 324 840
rect 336 828 348 840
rect 360 828 372 840
rect 384 828 396 840
rect 408 828 420 840
rect 432 828 444 840
rect 456 828 468 840
rect 480 828 492 840
rect 504 828 516 840
rect 528 828 540 840
rect 552 828 564 840
rect 576 828 588 840
rect 600 828 612 840
rect 624 828 636 840
rect 648 828 660 840
rect 672 828 684 840
rect 696 828 708 840
rect 720 828 732 840
rect 744 828 756 840
rect 768 828 780 840
rect 792 828 804 840
rect 816 828 828 840
rect 840 828 852 840
rect 864 828 876 840
rect 888 828 900 840
rect 912 828 924 840
rect 936 828 948 840
rect 960 828 972 840
rect 984 828 996 840
rect 1008 828 1020 840
rect 1032 828 1044 840
rect 1056 828 1068 840
rect 1080 828 1092 840
rect 1104 828 1116 840
rect 1128 828 1140 840
rect 1152 828 1164 840
rect 1176 828 1188 840
rect 1200 828 1212 840
rect 1224 828 1236 840
rect 1248 828 1260 840
rect 1272 828 1284 840
rect 1296 828 1308 840
rect 1320 828 1332 840
rect 1344 828 1356 840
rect 1368 828 1380 840
rect 1392 828 1404 840
rect 1416 828 1428 840
rect 1440 828 1452 840
rect 1464 828 1476 840
rect 1488 828 1500 840
rect 1512 828 1524 840
rect 1536 828 1548 840
rect 1560 828 1572 840
rect 1584 828 1596 840
rect 1608 828 1620 840
rect 1632 828 1644 840
rect 1656 828 1668 840
rect 1680 828 1692 840
rect 1704 828 1716 840
rect 1728 828 1740 840
rect 1752 828 1764 840
rect 1776 828 1788 840
rect 1800 828 1812 840
rect 1824 828 1836 840
rect 1848 828 1860 840
rect 1872 828 1884 840
rect 1896 828 1908 840
rect 1920 828 1932 840
rect 1944 828 1956 840
rect 1968 828 1980 840
rect 1992 828 2004 840
rect 2016 828 2028 840
rect 2040 828 2052 840
rect 2064 828 2076 840
rect 2088 828 2100 840
rect 2112 828 2124 840
rect 2136 828 2148 840
rect 2160 828 2172 840
rect 2184 828 2196 840
rect 2208 828 2220 840
rect 2232 828 2244 840
rect 2256 828 2268 840
rect 2280 828 2292 840
rect 2304 828 2316 840
rect 2328 828 2340 840
rect 2352 828 2364 840
rect 2376 828 2388 840
rect 2400 828 2412 840
rect 2424 828 2436 840
rect 2448 828 2460 840
rect 2472 828 2484 840
rect 2496 828 2508 840
rect 2520 828 2532 840
rect 2544 828 2556 840
rect 2568 828 2580 840
rect 2592 828 2604 840
rect 2616 828 2628 840
rect 2640 828 2652 840
rect 2664 828 2676 840
rect 2688 828 2700 840
rect 2712 828 2724 840
rect 2736 828 2748 840
rect 2760 828 2772 840
rect 2784 828 2796 840
rect 2808 828 2820 840
rect 2832 828 2844 840
rect 2856 828 2868 840
rect 2880 828 2892 840
rect 2904 828 2916 840
rect 2928 828 2940 840
rect 2952 828 2976 840
rect -1008 804 2976 828
rect -1008 792 -996 804
rect -984 792 -972 804
rect -960 792 -948 804
rect -936 792 -924 804
rect -912 792 -900 804
rect -888 792 -876 804
rect -864 792 -852 804
rect -840 792 -828 804
rect -816 792 -804 804
rect -792 792 -780 804
rect -768 792 -756 804
rect -744 792 -732 804
rect -720 792 -708 804
rect -696 792 -684 804
rect -672 792 -660 804
rect -648 792 -636 804
rect -624 792 -612 804
rect -600 792 -588 804
rect -576 792 -564 804
rect -552 792 -540 804
rect -528 792 -516 804
rect -504 792 -492 804
rect -480 792 -468 804
rect -456 792 -444 804
rect -432 792 -420 804
rect -408 792 -396 804
rect -384 792 -372 804
rect -360 792 -348 804
rect -336 792 -324 804
rect -312 792 -300 804
rect -288 792 -276 804
rect -264 792 -252 804
rect -240 792 -228 804
rect -216 792 -204 804
rect -192 792 -180 804
rect -168 792 -156 804
rect -144 792 -132 804
rect -120 792 -108 804
rect -96 792 -84 804
rect -72 792 -60 804
rect -48 792 -36 804
rect -24 792 -12 804
rect 0 792 12 804
rect 24 792 36 804
rect 48 792 60 804
rect 72 792 84 804
rect 96 792 108 804
rect 120 792 132 804
rect 144 792 156 804
rect 168 792 180 804
rect 192 792 204 804
rect 216 792 228 804
rect 240 792 252 804
rect 264 792 276 804
rect 288 792 300 804
rect 312 792 324 804
rect 336 792 348 804
rect 360 792 372 804
rect 384 792 396 804
rect 408 792 420 804
rect 432 792 444 804
rect 456 792 468 804
rect 480 792 492 804
rect 504 792 516 804
rect 528 792 540 804
rect 552 792 564 804
rect 576 792 588 804
rect 600 792 612 804
rect 624 792 636 804
rect 648 792 660 804
rect 672 792 684 804
rect 696 792 708 804
rect 720 792 732 804
rect 744 792 756 804
rect 768 792 780 804
rect 792 792 804 804
rect 816 792 828 804
rect 840 792 852 804
rect 864 792 876 804
rect 888 792 900 804
rect 912 792 924 804
rect 936 792 948 804
rect 960 792 972 804
rect 984 792 996 804
rect 1008 792 1020 804
rect 1032 792 1044 804
rect 1056 792 1068 804
rect 1080 792 1092 804
rect 1104 792 1116 804
rect 1128 792 1140 804
rect 1152 792 1164 804
rect 1176 792 1188 804
rect 1200 792 1212 804
rect 1224 792 1236 804
rect 1248 792 1260 804
rect 1272 792 1284 804
rect 1296 792 1308 804
rect 1320 792 1332 804
rect 1344 792 1356 804
rect 1368 792 1380 804
rect 1392 792 1404 804
rect 1416 792 1428 804
rect 1440 792 1452 804
rect 1464 792 1476 804
rect 1488 792 1500 804
rect 1512 792 1524 804
rect 1536 792 1548 804
rect 1560 792 1572 804
rect 1584 792 1596 804
rect 1608 792 1620 804
rect 1632 792 1644 804
rect 1656 792 1668 804
rect 1680 792 1692 804
rect 1704 792 1716 804
rect 1728 792 1740 804
rect 1752 792 1764 804
rect 1776 792 1788 804
rect 1800 792 1812 804
rect 1824 792 1836 804
rect 1848 792 1860 804
rect 1872 792 1884 804
rect 1896 792 1908 804
rect 1920 792 1932 804
rect 1944 792 1956 804
rect 1968 792 1980 804
rect 1992 792 2004 804
rect 2016 792 2028 804
rect 2040 792 2052 804
rect 2064 792 2076 804
rect 2088 792 2100 804
rect 2112 792 2124 804
rect 2136 792 2148 804
rect 2160 792 2172 804
rect 2184 792 2196 804
rect 2208 792 2220 804
rect 2232 792 2244 804
rect 2256 792 2268 804
rect 2280 792 2292 804
rect 2304 792 2316 804
rect 2328 792 2340 804
rect 2352 792 2364 804
rect 2376 792 2388 804
rect 2400 792 2412 804
rect 2424 792 2436 804
rect 2448 792 2460 804
rect 2472 792 2484 804
rect 2496 792 2508 804
rect 2520 792 2532 804
rect 2544 792 2556 804
rect 2568 792 2580 804
rect 2592 792 2604 804
rect 2616 792 2628 804
rect 2640 792 2652 804
rect 2664 792 2676 804
rect 2688 792 2700 804
rect 2712 792 2724 804
rect 2736 792 2748 804
rect 2760 792 2772 804
rect 2784 792 2796 804
rect 2808 792 2820 804
rect 2832 792 2844 804
rect 2856 792 2868 804
rect 2880 792 2892 804
rect 2904 792 2916 804
rect 2928 792 2940 804
rect 2952 792 2976 804
rect -1008 768 2976 792
rect -1008 756 -996 768
rect -984 756 -972 768
rect -960 756 -948 768
rect -936 756 -924 768
rect -912 756 -900 768
rect -888 756 -876 768
rect -864 756 -852 768
rect -840 756 -828 768
rect -816 756 -804 768
rect -792 756 -780 768
rect -768 756 -756 768
rect -744 756 -732 768
rect -720 756 -708 768
rect -696 756 -684 768
rect -672 756 -660 768
rect -648 756 -636 768
rect -624 756 -612 768
rect -600 756 -588 768
rect -576 756 -564 768
rect -552 756 -540 768
rect -528 756 -516 768
rect -504 756 -492 768
rect -480 756 -468 768
rect -456 756 -444 768
rect -432 756 -420 768
rect -408 756 -396 768
rect -384 756 -372 768
rect -360 756 -348 768
rect -336 756 -324 768
rect -312 756 -300 768
rect -288 756 -276 768
rect -264 756 -252 768
rect -240 756 -228 768
rect -216 756 -204 768
rect -192 756 -180 768
rect -168 756 -156 768
rect -144 756 -132 768
rect -120 756 -108 768
rect -96 756 -84 768
rect -72 756 -60 768
rect -48 756 -36 768
rect -24 756 -12 768
rect 0 756 12 768
rect 24 756 36 768
rect 48 756 60 768
rect 72 756 84 768
rect 96 756 108 768
rect 120 756 132 768
rect 144 756 156 768
rect 168 756 180 768
rect 192 756 204 768
rect 216 756 228 768
rect 240 756 252 768
rect 264 756 276 768
rect 288 756 300 768
rect 312 756 324 768
rect 336 756 348 768
rect 360 756 372 768
rect 384 756 396 768
rect 408 756 420 768
rect 432 756 444 768
rect 456 756 468 768
rect 480 756 492 768
rect 504 756 516 768
rect 528 756 540 768
rect 552 756 564 768
rect 576 756 588 768
rect 600 756 612 768
rect 624 756 636 768
rect 648 756 660 768
rect 672 756 684 768
rect 696 756 708 768
rect 720 756 732 768
rect 744 756 756 768
rect 768 756 780 768
rect 792 756 804 768
rect 816 756 828 768
rect 840 756 852 768
rect 864 756 876 768
rect 888 756 900 768
rect 912 756 924 768
rect 936 756 948 768
rect 960 756 972 768
rect 984 756 996 768
rect 1008 756 1020 768
rect 1032 756 1044 768
rect 1056 756 1068 768
rect 1080 756 1092 768
rect 1104 756 1116 768
rect 1128 756 1140 768
rect 1152 756 1164 768
rect 1176 756 1188 768
rect 1200 756 1212 768
rect 1224 756 1236 768
rect 1248 756 1260 768
rect 1272 756 1284 768
rect 1296 756 1308 768
rect 1320 756 1332 768
rect 1344 756 1356 768
rect 1368 756 1380 768
rect 1392 756 1404 768
rect 1416 756 1428 768
rect 1440 756 1452 768
rect 1464 756 1476 768
rect 1488 756 1500 768
rect 1512 756 1524 768
rect 1536 756 1548 768
rect 1560 756 1572 768
rect 1584 756 1596 768
rect 1608 756 1620 768
rect 1632 756 1644 768
rect 1656 756 1668 768
rect 1680 756 1692 768
rect 1704 756 1716 768
rect 1728 756 1740 768
rect 1752 756 1764 768
rect 1776 756 1788 768
rect 1800 756 1812 768
rect 1824 756 1836 768
rect 1848 756 1860 768
rect 1872 756 1884 768
rect 1896 756 1908 768
rect 1920 756 1932 768
rect 1944 756 1956 768
rect 1968 756 1980 768
rect 1992 756 2004 768
rect 2016 756 2028 768
rect 2040 756 2052 768
rect 2064 756 2076 768
rect 2088 756 2100 768
rect 2112 756 2124 768
rect 2136 756 2148 768
rect 2160 756 2172 768
rect 2184 756 2196 768
rect 2208 756 2220 768
rect 2232 756 2244 768
rect 2256 756 2268 768
rect 2280 756 2292 768
rect 2304 756 2316 768
rect 2328 756 2340 768
rect 2352 756 2364 768
rect 2376 756 2388 768
rect 2400 756 2412 768
rect 2424 756 2436 768
rect 2448 756 2460 768
rect 2472 756 2484 768
rect 2496 756 2508 768
rect 2520 756 2532 768
rect 2544 756 2556 768
rect 2568 756 2580 768
rect 2592 756 2604 768
rect 2616 756 2628 768
rect 2640 756 2652 768
rect 2664 756 2676 768
rect 2688 756 2700 768
rect 2712 756 2724 768
rect 2736 756 2748 768
rect 2760 756 2772 768
rect 2784 756 2796 768
rect 2808 756 2820 768
rect 2832 756 2844 768
rect 2856 756 2868 768
rect 2880 756 2892 768
rect 2904 756 2916 768
rect 2928 756 2940 768
rect 2952 756 2976 768
rect -1008 744 2976 756
rect -1008 -252 2976 -240
rect -1008 -264 -996 -252
rect -984 -264 -948 -252
rect -936 -264 -924 -252
rect -912 -264 -876 -252
rect -864 -264 -852 -252
rect -840 -264 -804 -252
rect -792 -264 -780 -252
rect -768 -264 -732 -252
rect -720 -264 -708 -252
rect -696 -264 -660 -252
rect -648 -264 -636 -252
rect -624 -264 -588 -252
rect -576 -264 -564 -252
rect -552 -264 -516 -252
rect -504 -264 -492 -252
rect -480 -264 -444 -252
rect -432 -264 -420 -252
rect -408 -264 -372 -252
rect -360 -264 -348 -252
rect -336 -264 -300 -252
rect -288 -264 -276 -252
rect -264 -264 -228 -252
rect -216 -264 -204 -252
rect -192 -264 -156 -252
rect -144 -264 -132 -252
rect -120 -264 -84 -252
rect -72 -264 -60 -252
rect -48 -264 -12 -252
rect 0 -264 12 -252
rect 24 -264 60 -252
rect 72 -264 84 -252
rect 96 -264 132 -252
rect 144 -264 156 -252
rect 168 -264 204 -252
rect 216 -264 228 -252
rect 240 -264 276 -252
rect 288 -264 300 -252
rect 312 -264 348 -252
rect 360 -264 372 -252
rect 384 -264 420 -252
rect 432 -264 444 -252
rect 456 -264 492 -252
rect 504 -264 516 -252
rect 528 -264 564 -252
rect 576 -264 588 -252
rect 600 -264 636 -252
rect 648 -264 660 -252
rect 672 -264 708 -252
rect 720 -264 732 -252
rect 744 -264 780 -252
rect 792 -264 804 -252
rect 816 -264 852 -252
rect 864 -264 876 -252
rect 888 -264 924 -252
rect 936 -264 948 -252
rect 960 -264 996 -252
rect 1008 -264 1020 -252
rect 1032 -264 1068 -252
rect 1080 -264 1092 -252
rect 1104 -264 1140 -252
rect 1152 -264 1164 -252
rect 1176 -264 1212 -252
rect 1224 -264 1236 -252
rect 1248 -264 1284 -252
rect 1296 -264 1308 -252
rect 1320 -264 1356 -252
rect 1368 -264 1380 -252
rect 1392 -264 1428 -252
rect 1440 -264 1452 -252
rect 1464 -264 1500 -252
rect 1512 -264 1524 -252
rect 1536 -264 1572 -252
rect 1584 -264 1596 -252
rect 1608 -264 1644 -252
rect 1656 -264 1668 -252
rect 1680 -264 1716 -252
rect 1728 -264 1740 -252
rect 1752 -264 1788 -252
rect 1800 -264 1812 -252
rect 1824 -264 1860 -252
rect 1872 -264 1884 -252
rect 1896 -264 1932 -252
rect 1944 -264 1956 -252
rect 1968 -264 2004 -252
rect 2016 -264 2028 -252
rect 2040 -264 2076 -252
rect 2088 -264 2100 -252
rect 2112 -264 2148 -252
rect 2160 -264 2172 -252
rect 2184 -264 2220 -252
rect 2232 -264 2244 -252
rect 2256 -264 2292 -252
rect 2304 -264 2316 -252
rect 2328 -264 2364 -252
rect 2376 -264 2388 -252
rect 2400 -264 2436 -252
rect 2448 -264 2460 -252
rect 2472 -264 2484 -252
rect 2496 -264 2532 -252
rect 2544 -264 2556 -252
rect 2568 -264 2604 -252
rect 2616 -264 2628 -252
rect 2640 -264 2676 -252
rect 2688 -264 2700 -252
rect 2712 -264 2724 -252
rect 2736 -264 2772 -252
rect 2784 -264 2796 -252
rect 2808 -264 2844 -252
rect 2856 -264 2868 -252
rect 2880 -264 2916 -252
rect 2928 -264 2940 -252
rect 2952 -264 2976 -252
rect -1008 -288 2976 -264
rect -1008 -300 -996 -288
rect -984 -300 -972 -288
rect -960 -300 -948 -288
rect -936 -300 -924 -288
rect -912 -300 -900 -288
rect -888 -300 -876 -288
rect -864 -300 -852 -288
rect -840 -300 -828 -288
rect -816 -300 -804 -288
rect -792 -300 -780 -288
rect -768 -300 -756 -288
rect -744 -300 -732 -288
rect -720 -300 -708 -288
rect -696 -300 -684 -288
rect -672 -300 -660 -288
rect -648 -300 -636 -288
rect -624 -300 -612 -288
rect -600 -300 -588 -288
rect -576 -300 -564 -288
rect -552 -300 -540 -288
rect -528 -300 -516 -288
rect -504 -300 -492 -288
rect -480 -300 -468 -288
rect -456 -300 -444 -288
rect -432 -300 -420 -288
rect -408 -300 -396 -288
rect -384 -300 -372 -288
rect -360 -300 -348 -288
rect -336 -300 -324 -288
rect -312 -300 -300 -288
rect -288 -300 -276 -288
rect -264 -300 -252 -288
rect -240 -300 -228 -288
rect -216 -300 -204 -288
rect -192 -300 -180 -288
rect -168 -300 -156 -288
rect -144 -300 -132 -288
rect -120 -300 -108 -288
rect -96 -300 -84 -288
rect -72 -300 -60 -288
rect -48 -300 -36 -288
rect -24 -300 -12 -288
rect 0 -300 12 -288
rect 24 -300 36 -288
rect 48 -300 60 -288
rect 72 -300 84 -288
rect 96 -300 108 -288
rect 120 -300 132 -288
rect 144 -300 156 -288
rect 168 -300 180 -288
rect 192 -300 204 -288
rect 216 -300 228 -288
rect 240 -300 252 -288
rect 264 -300 276 -288
rect 288 -300 300 -288
rect 312 -300 324 -288
rect 336 -300 348 -288
rect 360 -300 372 -288
rect 384 -300 396 -288
rect 408 -300 420 -288
rect 432 -300 444 -288
rect 456 -300 468 -288
rect 480 -300 492 -288
rect 504 -300 516 -288
rect 528 -300 540 -288
rect 552 -300 564 -288
rect 576 -300 588 -288
rect 600 -300 612 -288
rect 624 -300 636 -288
rect 648 -300 660 -288
rect 672 -300 684 -288
rect 696 -300 708 -288
rect 720 -300 732 -288
rect 744 -300 756 -288
rect 768 -300 780 -288
rect 792 -300 804 -288
rect 816 -300 828 -288
rect 840 -300 852 -288
rect 864 -300 876 -288
rect 888 -300 900 -288
rect 912 -300 924 -288
rect 936 -300 948 -288
rect 960 -300 972 -288
rect 984 -300 996 -288
rect 1008 -300 1020 -288
rect 1032 -300 1044 -288
rect 1056 -300 1068 -288
rect 1080 -300 1092 -288
rect 1104 -300 1116 -288
rect 1128 -300 1140 -288
rect 1152 -300 1164 -288
rect 1176 -300 1188 -288
rect 1200 -300 1212 -288
rect 1224 -300 1236 -288
rect 1248 -300 1260 -288
rect 1272 -300 1284 -288
rect 1296 -300 1308 -288
rect 1320 -300 1332 -288
rect 1344 -300 1356 -288
rect 1368 -300 1380 -288
rect 1392 -300 1404 -288
rect 1416 -300 1428 -288
rect 1440 -300 1452 -288
rect 1464 -300 1476 -288
rect 1488 -300 1500 -288
rect 1512 -300 1524 -288
rect 1536 -300 1548 -288
rect 1560 -300 1572 -288
rect 1584 -300 1596 -288
rect 1608 -300 1620 -288
rect 1632 -300 1644 -288
rect 1656 -300 1668 -288
rect 1680 -300 1692 -288
rect 1704 -300 1716 -288
rect 1728 -300 1740 -288
rect 1752 -300 1764 -288
rect 1776 -300 1788 -288
rect 1800 -300 1812 -288
rect 1824 -300 1836 -288
rect 1848 -300 1860 -288
rect 1872 -300 1884 -288
rect 1896 -300 1908 -288
rect 1920 -300 1932 -288
rect 1944 -300 1956 -288
rect 1968 -300 1980 -288
rect 1992 -300 2004 -288
rect 2016 -300 2028 -288
rect 2040 -300 2052 -288
rect 2064 -300 2076 -288
rect 2088 -300 2100 -288
rect 2112 -300 2124 -288
rect 2136 -300 2148 -288
rect 2160 -300 2172 -288
rect 2184 -300 2196 -288
rect 2208 -300 2220 -288
rect 2232 -300 2244 -288
rect 2256 -300 2268 -288
rect 2280 -300 2292 -288
rect 2304 -300 2316 -288
rect 2328 -300 2340 -288
rect 2352 -300 2364 -288
rect 2376 -300 2388 -288
rect 2400 -300 2412 -288
rect 2424 -300 2436 -288
rect 2448 -300 2460 -288
rect 2472 -300 2484 -288
rect 2496 -300 2508 -288
rect 2520 -300 2532 -288
rect 2544 -300 2556 -288
rect 2568 -300 2580 -288
rect 2592 -300 2604 -288
rect 2616 -300 2628 -288
rect 2640 -300 2652 -288
rect 2664 -300 2676 -288
rect 2688 -300 2700 -288
rect 2712 -300 2724 -288
rect 2736 -300 2748 -288
rect 2760 -300 2772 -288
rect 2784 -300 2796 -288
rect 2808 -300 2820 -288
rect 2832 -300 2844 -288
rect 2856 -300 2868 -288
rect 2880 -300 2892 -288
rect 2904 -300 2916 -288
rect 2928 -300 2940 -288
rect 2952 -300 2976 -288
rect -1008 -324 2976 -300
rect -1008 -336 -996 -324
rect -984 -336 -972 -324
rect -960 -336 -948 -324
rect -936 -336 -924 -324
rect -912 -336 -900 -324
rect -888 -336 -876 -324
rect -864 -336 -852 -324
rect -840 -336 -828 -324
rect -816 -336 -804 -324
rect -792 -336 -780 -324
rect -768 -336 -756 -324
rect -744 -336 -732 -324
rect -720 -336 -708 -324
rect -696 -336 -684 -324
rect -672 -336 -660 -324
rect -648 -336 -636 -324
rect -624 -336 -612 -324
rect -600 -336 -588 -324
rect -576 -336 -564 -324
rect -552 -336 -540 -324
rect -528 -336 -516 -324
rect -504 -336 -492 -324
rect -480 -336 -468 -324
rect -456 -336 -444 -324
rect -432 -336 -420 -324
rect -408 -336 -396 -324
rect -384 -336 -372 -324
rect -360 -336 -348 -324
rect -336 -336 -324 -324
rect -312 -336 -300 -324
rect -288 -336 -276 -324
rect -264 -336 -252 -324
rect -240 -336 -228 -324
rect -216 -336 -204 -324
rect -192 -336 -180 -324
rect -168 -336 -156 -324
rect -144 -336 -132 -324
rect -120 -336 -108 -324
rect -96 -336 -84 -324
rect -72 -336 -60 -324
rect -48 -336 -36 -324
rect -24 -336 -12 -324
rect 0 -336 12 -324
rect 24 -336 36 -324
rect 48 -336 60 -324
rect 72 -336 84 -324
rect 96 -336 108 -324
rect 120 -336 132 -324
rect 144 -336 156 -324
rect 168 -336 180 -324
rect 192 -336 204 -324
rect 216 -336 228 -324
rect 240 -336 252 -324
rect 264 -336 276 -324
rect 288 -336 300 -324
rect 312 -336 324 -324
rect 336 -336 348 -324
rect 360 -336 372 -324
rect 384 -336 396 -324
rect 408 -336 420 -324
rect 432 -336 444 -324
rect 456 -336 468 -324
rect 480 -336 492 -324
rect 504 -336 516 -324
rect 528 -336 540 -324
rect 552 -336 564 -324
rect 576 -336 588 -324
rect 600 -336 612 -324
rect 624 -336 636 -324
rect 648 -336 660 -324
rect 672 -336 684 -324
rect 696 -336 708 -324
rect 720 -336 732 -324
rect 744 -336 756 -324
rect 768 -336 780 -324
rect 792 -336 804 -324
rect 816 -336 828 -324
rect 840 -336 852 -324
rect 864 -336 876 -324
rect 888 -336 900 -324
rect 912 -336 924 -324
rect 936 -336 948 -324
rect 960 -336 972 -324
rect 984 -336 996 -324
rect 1008 -336 1020 -324
rect 1032 -336 1044 -324
rect 1056 -336 1068 -324
rect 1080 -336 1092 -324
rect 1104 -336 1116 -324
rect 1128 -336 1140 -324
rect 1152 -336 1164 -324
rect 1176 -336 1188 -324
rect 1200 -336 1212 -324
rect 1224 -336 1236 -324
rect 1248 -336 1260 -324
rect 1272 -336 1284 -324
rect 1296 -336 1308 -324
rect 1320 -336 1332 -324
rect 1344 -336 1356 -324
rect 1368 -336 1380 -324
rect 1392 -336 1404 -324
rect 1416 -336 1428 -324
rect 1440 -336 1452 -324
rect 1464 -336 1476 -324
rect 1488 -336 1500 -324
rect 1512 -336 1524 -324
rect 1536 -336 1548 -324
rect 1560 -336 1572 -324
rect 1584 -336 1596 -324
rect 1608 -336 1620 -324
rect 1632 -336 1644 -324
rect 1656 -336 1668 -324
rect 1680 -336 1692 -324
rect 1704 -336 1716 -324
rect 1728 -336 1740 -324
rect 1752 -336 1764 -324
rect 1776 -336 1788 -324
rect 1800 -336 1812 -324
rect 1824 -336 1836 -324
rect 1848 -336 1860 -324
rect 1872 -336 1884 -324
rect 1896 -336 1908 -324
rect 1920 -336 1932 -324
rect 1944 -336 1956 -324
rect 1968 -336 1980 -324
rect 1992 -336 2004 -324
rect 2016 -336 2028 -324
rect 2040 -336 2052 -324
rect 2064 -336 2076 -324
rect 2088 -336 2100 -324
rect 2112 -336 2124 -324
rect 2136 -336 2148 -324
rect 2160 -336 2172 -324
rect 2184 -336 2196 -324
rect 2208 -336 2220 -324
rect 2232 -336 2244 -324
rect 2256 -336 2268 -324
rect 2280 -336 2292 -324
rect 2304 -336 2316 -324
rect 2328 -336 2340 -324
rect 2352 -336 2364 -324
rect 2376 -336 2388 -324
rect 2400 -336 2412 -324
rect 2424 -336 2436 -324
rect 2448 -336 2460 -324
rect 2472 -336 2484 -324
rect 2496 -336 2508 -324
rect 2520 -336 2532 -324
rect 2544 -336 2556 -324
rect 2568 -336 2580 -324
rect 2592 -336 2604 -324
rect 2616 -336 2628 -324
rect 2640 -336 2652 -324
rect 2664 -336 2676 -324
rect 2688 -336 2700 -324
rect 2712 -336 2724 -324
rect 2736 -336 2748 -324
rect 2760 -336 2772 -324
rect 2784 -336 2796 -324
rect 2808 -336 2820 -324
rect 2832 -336 2844 -324
rect 2856 -336 2868 -324
rect 2880 -336 2892 -324
rect 2904 -336 2916 -324
rect 2928 -336 2940 -324
rect 2952 -336 2976 -324
rect -1008 -360 2976 -336
rect -1008 -372 -996 -360
rect -984 -372 -972 -360
rect -960 -372 -948 -360
rect -936 -372 -924 -360
rect -912 -372 -900 -360
rect -888 -372 -876 -360
rect -864 -372 -852 -360
rect -840 -372 -828 -360
rect -816 -372 -804 -360
rect -792 -372 -780 -360
rect -768 -372 -756 -360
rect -744 -372 -732 -360
rect -720 -372 -708 -360
rect -696 -372 -684 -360
rect -672 -372 -660 -360
rect -648 -372 -636 -360
rect -624 -372 -612 -360
rect -600 -372 -588 -360
rect -576 -372 -564 -360
rect -552 -372 -540 -360
rect -528 -372 -516 -360
rect -504 -372 -492 -360
rect -480 -372 -468 -360
rect -456 -372 -444 -360
rect -432 -372 -420 -360
rect -408 -372 -396 -360
rect -384 -372 -372 -360
rect -360 -372 -348 -360
rect -336 -372 -324 -360
rect -312 -372 -300 -360
rect -288 -372 -276 -360
rect -264 -372 -252 -360
rect -240 -372 -228 -360
rect -216 -372 -204 -360
rect -192 -372 -180 -360
rect -168 -372 -156 -360
rect -144 -372 -132 -360
rect -120 -372 -108 -360
rect -96 -372 -84 -360
rect -72 -372 -60 -360
rect -48 -372 -36 -360
rect -24 -372 -12 -360
rect 0 -372 12 -360
rect 24 -372 36 -360
rect 48 -372 60 -360
rect 72 -372 84 -360
rect 96 -372 108 -360
rect 120 -372 132 -360
rect 144 -372 156 -360
rect 168 -372 180 -360
rect 192 -372 204 -360
rect 216 -372 228 -360
rect 240 -372 252 -360
rect 264 -372 276 -360
rect 288 -372 300 -360
rect 312 -372 324 -360
rect 336 -372 348 -360
rect 360 -372 372 -360
rect 384 -372 396 -360
rect 408 -372 420 -360
rect 432 -372 444 -360
rect 456 -372 468 -360
rect 480 -372 492 -360
rect 504 -372 516 -360
rect 528 -372 540 -360
rect 552 -372 564 -360
rect 576 -372 588 -360
rect 600 -372 612 -360
rect 624 -372 636 -360
rect 648 -372 660 -360
rect 672 -372 684 -360
rect 696 -372 708 -360
rect 720 -372 732 -360
rect 744 -372 756 -360
rect 768 -372 780 -360
rect 792 -372 804 -360
rect 816 -372 828 -360
rect 840 -372 852 -360
rect 864 -372 876 -360
rect 888 -372 900 -360
rect 912 -372 924 -360
rect 936 -372 948 -360
rect 960 -372 972 -360
rect 984 -372 996 -360
rect 1008 -372 1020 -360
rect 1032 -372 1044 -360
rect 1056 -372 1068 -360
rect 1080 -372 1092 -360
rect 1104 -372 1116 -360
rect 1128 -372 1140 -360
rect 1152 -372 1164 -360
rect 1176 -372 1188 -360
rect 1200 -372 1212 -360
rect 1224 -372 1236 -360
rect 1248 -372 1260 -360
rect 1272 -372 1284 -360
rect 1296 -372 1308 -360
rect 1320 -372 1332 -360
rect 1344 -372 1356 -360
rect 1368 -372 1380 -360
rect 1392 -372 1404 -360
rect 1416 -372 1428 -360
rect 1440 -372 1452 -360
rect 1464 -372 1476 -360
rect 1488 -372 1500 -360
rect 1512 -372 1524 -360
rect 1536 -372 1548 -360
rect 1560 -372 1572 -360
rect 1584 -372 1596 -360
rect 1608 -372 1620 -360
rect 1632 -372 1644 -360
rect 1656 -372 1668 -360
rect 1680 -372 1692 -360
rect 1704 -372 1716 -360
rect 1728 -372 1740 -360
rect 1752 -372 1764 -360
rect 1776 -372 1788 -360
rect 1800 -372 1812 -360
rect 1824 -372 1836 -360
rect 1848 -372 1860 -360
rect 1872 -372 1884 -360
rect 1896 -372 1908 -360
rect 1920 -372 1932 -360
rect 1944 -372 1956 -360
rect 1968 -372 1980 -360
rect 1992 -372 2004 -360
rect 2016 -372 2028 -360
rect 2040 -372 2052 -360
rect 2064 -372 2076 -360
rect 2088 -372 2100 -360
rect 2112 -372 2124 -360
rect 2136 -372 2148 -360
rect 2160 -372 2172 -360
rect 2184 -372 2196 -360
rect 2208 -372 2220 -360
rect 2232 -372 2244 -360
rect 2256 -372 2268 -360
rect 2280 -372 2292 -360
rect 2304 -372 2316 -360
rect 2328 -372 2340 -360
rect 2352 -372 2364 -360
rect 2376 -372 2388 -360
rect 2400 -372 2412 -360
rect 2424 -372 2436 -360
rect 2448 -372 2460 -360
rect 2472 -372 2484 -360
rect 2496 -372 2508 -360
rect 2520 -372 2532 -360
rect 2544 -372 2556 -360
rect 2568 -372 2580 -360
rect 2592 -372 2604 -360
rect 2616 -372 2628 -360
rect 2640 -372 2652 -360
rect 2664 -372 2676 -360
rect 2688 -372 2700 -360
rect 2712 -372 2724 -360
rect 2736 -372 2748 -360
rect 2760 -372 2772 -360
rect 2784 -372 2796 -360
rect 2808 -372 2820 -360
rect 2832 -372 2844 -360
rect 2856 -372 2868 -360
rect 2880 -372 2892 -360
rect 2904 -372 2916 -360
rect 2928 -372 2940 -360
rect 2952 -372 2976 -360
rect -1008 -384 2976 -372
<< mimcapcontact >>
rect -996 864 -984 876
rect -948 864 -936 876
rect -924 864 -912 876
rect -876 864 -864 876
rect -852 864 -840 876
rect -804 864 -792 876
rect -780 864 -768 876
rect -732 864 -720 876
rect -708 864 -696 876
rect -660 864 -648 876
rect -636 864 -624 876
rect -588 864 -576 876
rect -564 864 -552 876
rect -516 864 -504 876
rect -492 864 -480 876
rect -444 864 -432 876
rect -420 864 -408 876
rect -372 864 -360 876
rect -348 864 -336 876
rect -300 864 -288 876
rect -276 864 -264 876
rect -228 864 -216 876
rect -204 864 -192 876
rect -156 864 -144 876
rect -132 864 -120 876
rect -84 864 -72 876
rect -60 864 -48 876
rect -12 864 0 876
rect 12 864 24 876
rect 60 864 72 876
rect 84 864 96 876
rect 132 864 144 876
rect 156 864 168 876
rect 204 864 216 876
rect 228 864 240 876
rect 276 864 288 876
rect 300 864 312 876
rect 348 864 360 876
rect 372 864 384 876
rect 420 864 432 876
rect 444 864 456 876
rect 492 864 504 876
rect 516 864 528 876
rect 564 864 576 876
rect 588 864 600 876
rect 636 864 648 876
rect 660 864 672 876
rect 708 864 720 876
rect 732 864 744 876
rect 780 864 792 876
rect 804 864 816 876
rect 852 864 864 876
rect 876 864 888 876
rect 924 864 936 876
rect 948 864 960 876
rect 996 864 1008 876
rect 1020 864 1032 876
rect 1068 864 1080 876
rect 1092 864 1104 876
rect 1140 864 1152 876
rect 1164 864 1176 876
rect 1212 864 1224 876
rect 1236 864 1248 876
rect 1284 864 1296 876
rect 1308 864 1320 876
rect 1356 864 1368 876
rect 1380 864 1392 876
rect 1428 864 1440 876
rect 1452 864 1464 876
rect 1500 864 1512 876
rect 1524 864 1536 876
rect 1572 864 1584 876
rect 1596 864 1608 876
rect 1644 864 1656 876
rect 1668 864 1680 876
rect 1716 864 1728 876
rect 1740 864 1752 876
rect 1788 864 1800 876
rect 1812 864 1824 876
rect 1860 864 1872 876
rect 1884 864 1896 876
rect 1932 864 1944 876
rect 1956 864 1968 876
rect 2004 864 2016 876
rect 2028 864 2040 876
rect 2076 864 2088 876
rect 2100 864 2112 876
rect 2148 864 2160 876
rect 2172 864 2184 876
rect 2220 864 2232 876
rect 2244 864 2256 876
rect 2292 864 2304 876
rect 2316 864 2328 876
rect 2364 864 2376 876
rect 2388 864 2400 876
rect 2436 864 2448 876
rect 2460 864 2472 876
rect 2484 864 2496 876
rect 2532 864 2544 876
rect 2556 864 2568 876
rect 2604 864 2616 876
rect 2628 864 2640 876
rect 2676 864 2688 876
rect 2700 864 2712 876
rect 2724 864 2736 876
rect 2772 864 2784 876
rect 2796 864 2808 876
rect 2844 864 2856 876
rect 2868 864 2880 876
rect 2916 864 2928 876
rect 2940 864 2952 876
rect -996 828 -984 840
rect -972 828 -960 840
rect -948 828 -936 840
rect -924 828 -912 840
rect -900 828 -888 840
rect -876 828 -864 840
rect -852 828 -840 840
rect -828 828 -816 840
rect -804 828 -792 840
rect -780 828 -768 840
rect -756 828 -744 840
rect -732 828 -720 840
rect -708 828 -696 840
rect -684 828 -672 840
rect -660 828 -648 840
rect -636 828 -624 840
rect -612 828 -600 840
rect -588 828 -576 840
rect -564 828 -552 840
rect -540 828 -528 840
rect -516 828 -504 840
rect -492 828 -480 840
rect -468 828 -456 840
rect -444 828 -432 840
rect -420 828 -408 840
rect -396 828 -384 840
rect -372 828 -360 840
rect -348 828 -336 840
rect -324 828 -312 840
rect -300 828 -288 840
rect -276 828 -264 840
rect -252 828 -240 840
rect -228 828 -216 840
rect -204 828 -192 840
rect -180 828 -168 840
rect -156 828 -144 840
rect -132 828 -120 840
rect -108 828 -96 840
rect -84 828 -72 840
rect -60 828 -48 840
rect -36 828 -24 840
rect -12 828 0 840
rect 12 828 24 840
rect 36 828 48 840
rect 60 828 72 840
rect 84 828 96 840
rect 108 828 120 840
rect 132 828 144 840
rect 156 828 168 840
rect 180 828 192 840
rect 204 828 216 840
rect 228 828 240 840
rect 252 828 264 840
rect 276 828 288 840
rect 300 828 312 840
rect 324 828 336 840
rect 348 828 360 840
rect 372 828 384 840
rect 396 828 408 840
rect 420 828 432 840
rect 444 828 456 840
rect 468 828 480 840
rect 492 828 504 840
rect 516 828 528 840
rect 540 828 552 840
rect 564 828 576 840
rect 588 828 600 840
rect 612 828 624 840
rect 636 828 648 840
rect 660 828 672 840
rect 684 828 696 840
rect 708 828 720 840
rect 732 828 744 840
rect 756 828 768 840
rect 780 828 792 840
rect 804 828 816 840
rect 828 828 840 840
rect 852 828 864 840
rect 876 828 888 840
rect 900 828 912 840
rect 924 828 936 840
rect 948 828 960 840
rect 972 828 984 840
rect 996 828 1008 840
rect 1020 828 1032 840
rect 1044 828 1056 840
rect 1068 828 1080 840
rect 1092 828 1104 840
rect 1116 828 1128 840
rect 1140 828 1152 840
rect 1164 828 1176 840
rect 1188 828 1200 840
rect 1212 828 1224 840
rect 1236 828 1248 840
rect 1260 828 1272 840
rect 1284 828 1296 840
rect 1308 828 1320 840
rect 1332 828 1344 840
rect 1356 828 1368 840
rect 1380 828 1392 840
rect 1404 828 1416 840
rect 1428 828 1440 840
rect 1452 828 1464 840
rect 1476 828 1488 840
rect 1500 828 1512 840
rect 1524 828 1536 840
rect 1548 828 1560 840
rect 1572 828 1584 840
rect 1596 828 1608 840
rect 1620 828 1632 840
rect 1644 828 1656 840
rect 1668 828 1680 840
rect 1692 828 1704 840
rect 1716 828 1728 840
rect 1740 828 1752 840
rect 1764 828 1776 840
rect 1788 828 1800 840
rect 1812 828 1824 840
rect 1836 828 1848 840
rect 1860 828 1872 840
rect 1884 828 1896 840
rect 1908 828 1920 840
rect 1932 828 1944 840
rect 1956 828 1968 840
rect 1980 828 1992 840
rect 2004 828 2016 840
rect 2028 828 2040 840
rect 2052 828 2064 840
rect 2076 828 2088 840
rect 2100 828 2112 840
rect 2124 828 2136 840
rect 2148 828 2160 840
rect 2172 828 2184 840
rect 2196 828 2208 840
rect 2220 828 2232 840
rect 2244 828 2256 840
rect 2268 828 2280 840
rect 2292 828 2304 840
rect 2316 828 2328 840
rect 2340 828 2352 840
rect 2364 828 2376 840
rect 2388 828 2400 840
rect 2412 828 2424 840
rect 2436 828 2448 840
rect 2460 828 2472 840
rect 2484 828 2496 840
rect 2508 828 2520 840
rect 2532 828 2544 840
rect 2556 828 2568 840
rect 2580 828 2592 840
rect 2604 828 2616 840
rect 2628 828 2640 840
rect 2652 828 2664 840
rect 2676 828 2688 840
rect 2700 828 2712 840
rect 2724 828 2736 840
rect 2748 828 2760 840
rect 2772 828 2784 840
rect 2796 828 2808 840
rect 2820 828 2832 840
rect 2844 828 2856 840
rect 2868 828 2880 840
rect 2892 828 2904 840
rect 2916 828 2928 840
rect 2940 828 2952 840
rect -996 792 -984 804
rect -972 792 -960 804
rect -948 792 -936 804
rect -924 792 -912 804
rect -900 792 -888 804
rect -876 792 -864 804
rect -852 792 -840 804
rect -828 792 -816 804
rect -804 792 -792 804
rect -780 792 -768 804
rect -756 792 -744 804
rect -732 792 -720 804
rect -708 792 -696 804
rect -684 792 -672 804
rect -660 792 -648 804
rect -636 792 -624 804
rect -612 792 -600 804
rect -588 792 -576 804
rect -564 792 -552 804
rect -540 792 -528 804
rect -516 792 -504 804
rect -492 792 -480 804
rect -468 792 -456 804
rect -444 792 -432 804
rect -420 792 -408 804
rect -396 792 -384 804
rect -372 792 -360 804
rect -348 792 -336 804
rect -324 792 -312 804
rect -300 792 -288 804
rect -276 792 -264 804
rect -252 792 -240 804
rect -228 792 -216 804
rect -204 792 -192 804
rect -180 792 -168 804
rect -156 792 -144 804
rect -132 792 -120 804
rect -108 792 -96 804
rect -84 792 -72 804
rect -60 792 -48 804
rect -36 792 -24 804
rect -12 792 0 804
rect 12 792 24 804
rect 36 792 48 804
rect 60 792 72 804
rect 84 792 96 804
rect 108 792 120 804
rect 132 792 144 804
rect 156 792 168 804
rect 180 792 192 804
rect 204 792 216 804
rect 228 792 240 804
rect 252 792 264 804
rect 276 792 288 804
rect 300 792 312 804
rect 324 792 336 804
rect 348 792 360 804
rect 372 792 384 804
rect 396 792 408 804
rect 420 792 432 804
rect 444 792 456 804
rect 468 792 480 804
rect 492 792 504 804
rect 516 792 528 804
rect 540 792 552 804
rect 564 792 576 804
rect 588 792 600 804
rect 612 792 624 804
rect 636 792 648 804
rect 660 792 672 804
rect 684 792 696 804
rect 708 792 720 804
rect 732 792 744 804
rect 756 792 768 804
rect 780 792 792 804
rect 804 792 816 804
rect 828 792 840 804
rect 852 792 864 804
rect 876 792 888 804
rect 900 792 912 804
rect 924 792 936 804
rect 948 792 960 804
rect 972 792 984 804
rect 996 792 1008 804
rect 1020 792 1032 804
rect 1044 792 1056 804
rect 1068 792 1080 804
rect 1092 792 1104 804
rect 1116 792 1128 804
rect 1140 792 1152 804
rect 1164 792 1176 804
rect 1188 792 1200 804
rect 1212 792 1224 804
rect 1236 792 1248 804
rect 1260 792 1272 804
rect 1284 792 1296 804
rect 1308 792 1320 804
rect 1332 792 1344 804
rect 1356 792 1368 804
rect 1380 792 1392 804
rect 1404 792 1416 804
rect 1428 792 1440 804
rect 1452 792 1464 804
rect 1476 792 1488 804
rect 1500 792 1512 804
rect 1524 792 1536 804
rect 1548 792 1560 804
rect 1572 792 1584 804
rect 1596 792 1608 804
rect 1620 792 1632 804
rect 1644 792 1656 804
rect 1668 792 1680 804
rect 1692 792 1704 804
rect 1716 792 1728 804
rect 1740 792 1752 804
rect 1764 792 1776 804
rect 1788 792 1800 804
rect 1812 792 1824 804
rect 1836 792 1848 804
rect 1860 792 1872 804
rect 1884 792 1896 804
rect 1908 792 1920 804
rect 1932 792 1944 804
rect 1956 792 1968 804
rect 1980 792 1992 804
rect 2004 792 2016 804
rect 2028 792 2040 804
rect 2052 792 2064 804
rect 2076 792 2088 804
rect 2100 792 2112 804
rect 2124 792 2136 804
rect 2148 792 2160 804
rect 2172 792 2184 804
rect 2196 792 2208 804
rect 2220 792 2232 804
rect 2244 792 2256 804
rect 2268 792 2280 804
rect 2292 792 2304 804
rect 2316 792 2328 804
rect 2340 792 2352 804
rect 2364 792 2376 804
rect 2388 792 2400 804
rect 2412 792 2424 804
rect 2436 792 2448 804
rect 2460 792 2472 804
rect 2484 792 2496 804
rect 2508 792 2520 804
rect 2532 792 2544 804
rect 2556 792 2568 804
rect 2580 792 2592 804
rect 2604 792 2616 804
rect 2628 792 2640 804
rect 2652 792 2664 804
rect 2676 792 2688 804
rect 2700 792 2712 804
rect 2724 792 2736 804
rect 2748 792 2760 804
rect 2772 792 2784 804
rect 2796 792 2808 804
rect 2820 792 2832 804
rect 2844 792 2856 804
rect 2868 792 2880 804
rect 2892 792 2904 804
rect 2916 792 2928 804
rect 2940 792 2952 804
rect -996 756 -984 768
rect -972 756 -960 768
rect -948 756 -936 768
rect -924 756 -912 768
rect -900 756 -888 768
rect -876 756 -864 768
rect -852 756 -840 768
rect -828 756 -816 768
rect -804 756 -792 768
rect -780 756 -768 768
rect -756 756 -744 768
rect -732 756 -720 768
rect -708 756 -696 768
rect -684 756 -672 768
rect -660 756 -648 768
rect -636 756 -624 768
rect -612 756 -600 768
rect -588 756 -576 768
rect -564 756 -552 768
rect -540 756 -528 768
rect -516 756 -504 768
rect -492 756 -480 768
rect -468 756 -456 768
rect -444 756 -432 768
rect -420 756 -408 768
rect -396 756 -384 768
rect -372 756 -360 768
rect -348 756 -336 768
rect -324 756 -312 768
rect -300 756 -288 768
rect -276 756 -264 768
rect -252 756 -240 768
rect -228 756 -216 768
rect -204 756 -192 768
rect -180 756 -168 768
rect -156 756 -144 768
rect -132 756 -120 768
rect -108 756 -96 768
rect -84 756 -72 768
rect -60 756 -48 768
rect -36 756 -24 768
rect -12 756 0 768
rect 12 756 24 768
rect 36 756 48 768
rect 60 756 72 768
rect 84 756 96 768
rect 108 756 120 768
rect 132 756 144 768
rect 156 756 168 768
rect 180 756 192 768
rect 204 756 216 768
rect 228 756 240 768
rect 252 756 264 768
rect 276 756 288 768
rect 300 756 312 768
rect 324 756 336 768
rect 348 756 360 768
rect 372 756 384 768
rect 396 756 408 768
rect 420 756 432 768
rect 444 756 456 768
rect 468 756 480 768
rect 492 756 504 768
rect 516 756 528 768
rect 540 756 552 768
rect 564 756 576 768
rect 588 756 600 768
rect 612 756 624 768
rect 636 756 648 768
rect 660 756 672 768
rect 684 756 696 768
rect 708 756 720 768
rect 732 756 744 768
rect 756 756 768 768
rect 780 756 792 768
rect 804 756 816 768
rect 828 756 840 768
rect 852 756 864 768
rect 876 756 888 768
rect 900 756 912 768
rect 924 756 936 768
rect 948 756 960 768
rect 972 756 984 768
rect 996 756 1008 768
rect 1020 756 1032 768
rect 1044 756 1056 768
rect 1068 756 1080 768
rect 1092 756 1104 768
rect 1116 756 1128 768
rect 1140 756 1152 768
rect 1164 756 1176 768
rect 1188 756 1200 768
rect 1212 756 1224 768
rect 1236 756 1248 768
rect 1260 756 1272 768
rect 1284 756 1296 768
rect 1308 756 1320 768
rect 1332 756 1344 768
rect 1356 756 1368 768
rect 1380 756 1392 768
rect 1404 756 1416 768
rect 1428 756 1440 768
rect 1452 756 1464 768
rect 1476 756 1488 768
rect 1500 756 1512 768
rect 1524 756 1536 768
rect 1548 756 1560 768
rect 1572 756 1584 768
rect 1596 756 1608 768
rect 1620 756 1632 768
rect 1644 756 1656 768
rect 1668 756 1680 768
rect 1692 756 1704 768
rect 1716 756 1728 768
rect 1740 756 1752 768
rect 1764 756 1776 768
rect 1788 756 1800 768
rect 1812 756 1824 768
rect 1836 756 1848 768
rect 1860 756 1872 768
rect 1884 756 1896 768
rect 1908 756 1920 768
rect 1932 756 1944 768
rect 1956 756 1968 768
rect 1980 756 1992 768
rect 2004 756 2016 768
rect 2028 756 2040 768
rect 2052 756 2064 768
rect 2076 756 2088 768
rect 2100 756 2112 768
rect 2124 756 2136 768
rect 2148 756 2160 768
rect 2172 756 2184 768
rect 2196 756 2208 768
rect 2220 756 2232 768
rect 2244 756 2256 768
rect 2268 756 2280 768
rect 2292 756 2304 768
rect 2316 756 2328 768
rect 2340 756 2352 768
rect 2364 756 2376 768
rect 2388 756 2400 768
rect 2412 756 2424 768
rect 2436 756 2448 768
rect 2460 756 2472 768
rect 2484 756 2496 768
rect 2508 756 2520 768
rect 2532 756 2544 768
rect 2556 756 2568 768
rect 2580 756 2592 768
rect 2604 756 2616 768
rect 2628 756 2640 768
rect 2652 756 2664 768
rect 2676 756 2688 768
rect 2700 756 2712 768
rect 2724 756 2736 768
rect 2748 756 2760 768
rect 2772 756 2784 768
rect 2796 756 2808 768
rect 2820 756 2832 768
rect 2844 756 2856 768
rect 2868 756 2880 768
rect 2892 756 2904 768
rect 2916 756 2928 768
rect 2940 756 2952 768
rect -996 -264 -984 -252
rect -948 -264 -936 -252
rect -924 -264 -912 -252
rect -876 -264 -864 -252
rect -852 -264 -840 -252
rect -804 -264 -792 -252
rect -780 -264 -768 -252
rect -732 -264 -720 -252
rect -708 -264 -696 -252
rect -660 -264 -648 -252
rect -636 -264 -624 -252
rect -588 -264 -576 -252
rect -564 -264 -552 -252
rect -516 -264 -504 -252
rect -492 -264 -480 -252
rect -444 -264 -432 -252
rect -420 -264 -408 -252
rect -372 -264 -360 -252
rect -348 -264 -336 -252
rect -300 -264 -288 -252
rect -276 -264 -264 -252
rect -228 -264 -216 -252
rect -204 -264 -192 -252
rect -156 -264 -144 -252
rect -132 -264 -120 -252
rect -84 -264 -72 -252
rect -60 -264 -48 -252
rect -12 -264 0 -252
rect 12 -264 24 -252
rect 60 -264 72 -252
rect 84 -264 96 -252
rect 132 -264 144 -252
rect 156 -264 168 -252
rect 204 -264 216 -252
rect 228 -264 240 -252
rect 276 -264 288 -252
rect 300 -264 312 -252
rect 348 -264 360 -252
rect 372 -264 384 -252
rect 420 -264 432 -252
rect 444 -264 456 -252
rect 492 -264 504 -252
rect 516 -264 528 -252
rect 564 -264 576 -252
rect 588 -264 600 -252
rect 636 -264 648 -252
rect 660 -264 672 -252
rect 708 -264 720 -252
rect 732 -264 744 -252
rect 780 -264 792 -252
rect 804 -264 816 -252
rect 852 -264 864 -252
rect 876 -264 888 -252
rect 924 -264 936 -252
rect 948 -264 960 -252
rect 996 -264 1008 -252
rect 1020 -264 1032 -252
rect 1068 -264 1080 -252
rect 1092 -264 1104 -252
rect 1140 -264 1152 -252
rect 1164 -264 1176 -252
rect 1212 -264 1224 -252
rect 1236 -264 1248 -252
rect 1284 -264 1296 -252
rect 1308 -264 1320 -252
rect 1356 -264 1368 -252
rect 1380 -264 1392 -252
rect 1428 -264 1440 -252
rect 1452 -264 1464 -252
rect 1500 -264 1512 -252
rect 1524 -264 1536 -252
rect 1572 -264 1584 -252
rect 1596 -264 1608 -252
rect 1644 -264 1656 -252
rect 1668 -264 1680 -252
rect 1716 -264 1728 -252
rect 1740 -264 1752 -252
rect 1788 -264 1800 -252
rect 1812 -264 1824 -252
rect 1860 -264 1872 -252
rect 1884 -264 1896 -252
rect 1932 -264 1944 -252
rect 1956 -264 1968 -252
rect 2004 -264 2016 -252
rect 2028 -264 2040 -252
rect 2076 -264 2088 -252
rect 2100 -264 2112 -252
rect 2148 -264 2160 -252
rect 2172 -264 2184 -252
rect 2220 -264 2232 -252
rect 2244 -264 2256 -252
rect 2292 -264 2304 -252
rect 2316 -264 2328 -252
rect 2364 -264 2376 -252
rect 2388 -264 2400 -252
rect 2436 -264 2448 -252
rect 2460 -264 2472 -252
rect 2484 -264 2496 -252
rect 2532 -264 2544 -252
rect 2556 -264 2568 -252
rect 2604 -264 2616 -252
rect 2628 -264 2640 -252
rect 2676 -264 2688 -252
rect 2700 -264 2712 -252
rect 2724 -264 2736 -252
rect 2772 -264 2784 -252
rect 2796 -264 2808 -252
rect 2844 -264 2856 -252
rect 2868 -264 2880 -252
rect 2916 -264 2928 -252
rect 2940 -264 2952 -252
rect -996 -300 -984 -288
rect -972 -300 -960 -288
rect -948 -300 -936 -288
rect -924 -300 -912 -288
rect -900 -300 -888 -288
rect -876 -300 -864 -288
rect -852 -300 -840 -288
rect -828 -300 -816 -288
rect -804 -300 -792 -288
rect -780 -300 -768 -288
rect -756 -300 -744 -288
rect -732 -300 -720 -288
rect -708 -300 -696 -288
rect -684 -300 -672 -288
rect -660 -300 -648 -288
rect -636 -300 -624 -288
rect -612 -300 -600 -288
rect -588 -300 -576 -288
rect -564 -300 -552 -288
rect -540 -300 -528 -288
rect -516 -300 -504 -288
rect -492 -300 -480 -288
rect -468 -300 -456 -288
rect -444 -300 -432 -288
rect -420 -300 -408 -288
rect -396 -300 -384 -288
rect -372 -300 -360 -288
rect -348 -300 -336 -288
rect -324 -300 -312 -288
rect -300 -300 -288 -288
rect -276 -300 -264 -288
rect -252 -300 -240 -288
rect -228 -300 -216 -288
rect -204 -300 -192 -288
rect -180 -300 -168 -288
rect -156 -300 -144 -288
rect -132 -300 -120 -288
rect -108 -300 -96 -288
rect -84 -300 -72 -288
rect -60 -300 -48 -288
rect -36 -300 -24 -288
rect -12 -300 0 -288
rect 12 -300 24 -288
rect 36 -300 48 -288
rect 60 -300 72 -288
rect 84 -300 96 -288
rect 108 -300 120 -288
rect 132 -300 144 -288
rect 156 -300 168 -288
rect 180 -300 192 -288
rect 204 -300 216 -288
rect 228 -300 240 -288
rect 252 -300 264 -288
rect 276 -300 288 -288
rect 300 -300 312 -288
rect 324 -300 336 -288
rect 348 -300 360 -288
rect 372 -300 384 -288
rect 396 -300 408 -288
rect 420 -300 432 -288
rect 444 -300 456 -288
rect 468 -300 480 -288
rect 492 -300 504 -288
rect 516 -300 528 -288
rect 540 -300 552 -288
rect 564 -300 576 -288
rect 588 -300 600 -288
rect 612 -300 624 -288
rect 636 -300 648 -288
rect 660 -300 672 -288
rect 684 -300 696 -288
rect 708 -300 720 -288
rect 732 -300 744 -288
rect 756 -300 768 -288
rect 780 -300 792 -288
rect 804 -300 816 -288
rect 828 -300 840 -288
rect 852 -300 864 -288
rect 876 -300 888 -288
rect 900 -300 912 -288
rect 924 -300 936 -288
rect 948 -300 960 -288
rect 972 -300 984 -288
rect 996 -300 1008 -288
rect 1020 -300 1032 -288
rect 1044 -300 1056 -288
rect 1068 -300 1080 -288
rect 1092 -300 1104 -288
rect 1116 -300 1128 -288
rect 1140 -300 1152 -288
rect 1164 -300 1176 -288
rect 1188 -300 1200 -288
rect 1212 -300 1224 -288
rect 1236 -300 1248 -288
rect 1260 -300 1272 -288
rect 1284 -300 1296 -288
rect 1308 -300 1320 -288
rect 1332 -300 1344 -288
rect 1356 -300 1368 -288
rect 1380 -300 1392 -288
rect 1404 -300 1416 -288
rect 1428 -300 1440 -288
rect 1452 -300 1464 -288
rect 1476 -300 1488 -288
rect 1500 -300 1512 -288
rect 1524 -300 1536 -288
rect 1548 -300 1560 -288
rect 1572 -300 1584 -288
rect 1596 -300 1608 -288
rect 1620 -300 1632 -288
rect 1644 -300 1656 -288
rect 1668 -300 1680 -288
rect 1692 -300 1704 -288
rect 1716 -300 1728 -288
rect 1740 -300 1752 -288
rect 1764 -300 1776 -288
rect 1788 -300 1800 -288
rect 1812 -300 1824 -288
rect 1836 -300 1848 -288
rect 1860 -300 1872 -288
rect 1884 -300 1896 -288
rect 1908 -300 1920 -288
rect 1932 -300 1944 -288
rect 1956 -300 1968 -288
rect 1980 -300 1992 -288
rect 2004 -300 2016 -288
rect 2028 -300 2040 -288
rect 2052 -300 2064 -288
rect 2076 -300 2088 -288
rect 2100 -300 2112 -288
rect 2124 -300 2136 -288
rect 2148 -300 2160 -288
rect 2172 -300 2184 -288
rect 2196 -300 2208 -288
rect 2220 -300 2232 -288
rect 2244 -300 2256 -288
rect 2268 -300 2280 -288
rect 2292 -300 2304 -288
rect 2316 -300 2328 -288
rect 2340 -300 2352 -288
rect 2364 -300 2376 -288
rect 2388 -300 2400 -288
rect 2412 -300 2424 -288
rect 2436 -300 2448 -288
rect 2460 -300 2472 -288
rect 2484 -300 2496 -288
rect 2508 -300 2520 -288
rect 2532 -300 2544 -288
rect 2556 -300 2568 -288
rect 2580 -300 2592 -288
rect 2604 -300 2616 -288
rect 2628 -300 2640 -288
rect 2652 -300 2664 -288
rect 2676 -300 2688 -288
rect 2700 -300 2712 -288
rect 2724 -300 2736 -288
rect 2748 -300 2760 -288
rect 2772 -300 2784 -288
rect 2796 -300 2808 -288
rect 2820 -300 2832 -288
rect 2844 -300 2856 -288
rect 2868 -300 2880 -288
rect 2892 -300 2904 -288
rect 2916 -300 2928 -288
rect 2940 -300 2952 -288
rect -996 -336 -984 -324
rect -972 -336 -960 -324
rect -948 -336 -936 -324
rect -924 -336 -912 -324
rect -900 -336 -888 -324
rect -876 -336 -864 -324
rect -852 -336 -840 -324
rect -828 -336 -816 -324
rect -804 -336 -792 -324
rect -780 -336 -768 -324
rect -756 -336 -744 -324
rect -732 -336 -720 -324
rect -708 -336 -696 -324
rect -684 -336 -672 -324
rect -660 -336 -648 -324
rect -636 -336 -624 -324
rect -612 -336 -600 -324
rect -588 -336 -576 -324
rect -564 -336 -552 -324
rect -540 -336 -528 -324
rect -516 -336 -504 -324
rect -492 -336 -480 -324
rect -468 -336 -456 -324
rect -444 -336 -432 -324
rect -420 -336 -408 -324
rect -396 -336 -384 -324
rect -372 -336 -360 -324
rect -348 -336 -336 -324
rect -324 -336 -312 -324
rect -300 -336 -288 -324
rect -276 -336 -264 -324
rect -252 -336 -240 -324
rect -228 -336 -216 -324
rect -204 -336 -192 -324
rect -180 -336 -168 -324
rect -156 -336 -144 -324
rect -132 -336 -120 -324
rect -108 -336 -96 -324
rect -84 -336 -72 -324
rect -60 -336 -48 -324
rect -36 -336 -24 -324
rect -12 -336 0 -324
rect 12 -336 24 -324
rect 36 -336 48 -324
rect 60 -336 72 -324
rect 84 -336 96 -324
rect 108 -336 120 -324
rect 132 -336 144 -324
rect 156 -336 168 -324
rect 180 -336 192 -324
rect 204 -336 216 -324
rect 228 -336 240 -324
rect 252 -336 264 -324
rect 276 -336 288 -324
rect 300 -336 312 -324
rect 324 -336 336 -324
rect 348 -336 360 -324
rect 372 -336 384 -324
rect 396 -336 408 -324
rect 420 -336 432 -324
rect 444 -336 456 -324
rect 468 -336 480 -324
rect 492 -336 504 -324
rect 516 -336 528 -324
rect 540 -336 552 -324
rect 564 -336 576 -324
rect 588 -336 600 -324
rect 612 -336 624 -324
rect 636 -336 648 -324
rect 660 -336 672 -324
rect 684 -336 696 -324
rect 708 -336 720 -324
rect 732 -336 744 -324
rect 756 -336 768 -324
rect 780 -336 792 -324
rect 804 -336 816 -324
rect 828 -336 840 -324
rect 852 -336 864 -324
rect 876 -336 888 -324
rect 900 -336 912 -324
rect 924 -336 936 -324
rect 948 -336 960 -324
rect 972 -336 984 -324
rect 996 -336 1008 -324
rect 1020 -336 1032 -324
rect 1044 -336 1056 -324
rect 1068 -336 1080 -324
rect 1092 -336 1104 -324
rect 1116 -336 1128 -324
rect 1140 -336 1152 -324
rect 1164 -336 1176 -324
rect 1188 -336 1200 -324
rect 1212 -336 1224 -324
rect 1236 -336 1248 -324
rect 1260 -336 1272 -324
rect 1284 -336 1296 -324
rect 1308 -336 1320 -324
rect 1332 -336 1344 -324
rect 1356 -336 1368 -324
rect 1380 -336 1392 -324
rect 1404 -336 1416 -324
rect 1428 -336 1440 -324
rect 1452 -336 1464 -324
rect 1476 -336 1488 -324
rect 1500 -336 1512 -324
rect 1524 -336 1536 -324
rect 1548 -336 1560 -324
rect 1572 -336 1584 -324
rect 1596 -336 1608 -324
rect 1620 -336 1632 -324
rect 1644 -336 1656 -324
rect 1668 -336 1680 -324
rect 1692 -336 1704 -324
rect 1716 -336 1728 -324
rect 1740 -336 1752 -324
rect 1764 -336 1776 -324
rect 1788 -336 1800 -324
rect 1812 -336 1824 -324
rect 1836 -336 1848 -324
rect 1860 -336 1872 -324
rect 1884 -336 1896 -324
rect 1908 -336 1920 -324
rect 1932 -336 1944 -324
rect 1956 -336 1968 -324
rect 1980 -336 1992 -324
rect 2004 -336 2016 -324
rect 2028 -336 2040 -324
rect 2052 -336 2064 -324
rect 2076 -336 2088 -324
rect 2100 -336 2112 -324
rect 2124 -336 2136 -324
rect 2148 -336 2160 -324
rect 2172 -336 2184 -324
rect 2196 -336 2208 -324
rect 2220 -336 2232 -324
rect 2244 -336 2256 -324
rect 2268 -336 2280 -324
rect 2292 -336 2304 -324
rect 2316 -336 2328 -324
rect 2340 -336 2352 -324
rect 2364 -336 2376 -324
rect 2388 -336 2400 -324
rect 2412 -336 2424 -324
rect 2436 -336 2448 -324
rect 2460 -336 2472 -324
rect 2484 -336 2496 -324
rect 2508 -336 2520 -324
rect 2532 -336 2544 -324
rect 2556 -336 2568 -324
rect 2580 -336 2592 -324
rect 2604 -336 2616 -324
rect 2628 -336 2640 -324
rect 2652 -336 2664 -324
rect 2676 -336 2688 -324
rect 2700 -336 2712 -324
rect 2724 -336 2736 -324
rect 2748 -336 2760 -324
rect 2772 -336 2784 -324
rect 2796 -336 2808 -324
rect 2820 -336 2832 -324
rect 2844 -336 2856 -324
rect 2868 -336 2880 -324
rect 2892 -336 2904 -324
rect 2916 -336 2928 -324
rect 2940 -336 2952 -324
rect -996 -372 -984 -360
rect -972 -372 -960 -360
rect -948 -372 -936 -360
rect -924 -372 -912 -360
rect -900 -372 -888 -360
rect -876 -372 -864 -360
rect -852 -372 -840 -360
rect -828 -372 -816 -360
rect -804 -372 -792 -360
rect -780 -372 -768 -360
rect -756 -372 -744 -360
rect -732 -372 -720 -360
rect -708 -372 -696 -360
rect -684 -372 -672 -360
rect -660 -372 -648 -360
rect -636 -372 -624 -360
rect -612 -372 -600 -360
rect -588 -372 -576 -360
rect -564 -372 -552 -360
rect -540 -372 -528 -360
rect -516 -372 -504 -360
rect -492 -372 -480 -360
rect -468 -372 -456 -360
rect -444 -372 -432 -360
rect -420 -372 -408 -360
rect -396 -372 -384 -360
rect -372 -372 -360 -360
rect -348 -372 -336 -360
rect -324 -372 -312 -360
rect -300 -372 -288 -360
rect -276 -372 -264 -360
rect -252 -372 -240 -360
rect -228 -372 -216 -360
rect -204 -372 -192 -360
rect -180 -372 -168 -360
rect -156 -372 -144 -360
rect -132 -372 -120 -360
rect -108 -372 -96 -360
rect -84 -372 -72 -360
rect -60 -372 -48 -360
rect -36 -372 -24 -360
rect -12 -372 0 -360
rect 12 -372 24 -360
rect 36 -372 48 -360
rect 60 -372 72 -360
rect 84 -372 96 -360
rect 108 -372 120 -360
rect 132 -372 144 -360
rect 156 -372 168 -360
rect 180 -372 192 -360
rect 204 -372 216 -360
rect 228 -372 240 -360
rect 252 -372 264 -360
rect 276 -372 288 -360
rect 300 -372 312 -360
rect 324 -372 336 -360
rect 348 -372 360 -360
rect 372 -372 384 -360
rect 396 -372 408 -360
rect 420 -372 432 -360
rect 444 -372 456 -360
rect 468 -372 480 -360
rect 492 -372 504 -360
rect 516 -372 528 -360
rect 540 -372 552 -360
rect 564 -372 576 -360
rect 588 -372 600 -360
rect 612 -372 624 -360
rect 636 -372 648 -360
rect 660 -372 672 -360
rect 684 -372 696 -360
rect 708 -372 720 -360
rect 732 -372 744 -360
rect 756 -372 768 -360
rect 780 -372 792 -360
rect 804 -372 816 -360
rect 828 -372 840 -360
rect 852 -372 864 -360
rect 876 -372 888 -360
rect 900 -372 912 -360
rect 924 -372 936 -360
rect 948 -372 960 -360
rect 972 -372 984 -360
rect 996 -372 1008 -360
rect 1020 -372 1032 -360
rect 1044 -372 1056 -360
rect 1068 -372 1080 -360
rect 1092 -372 1104 -360
rect 1116 -372 1128 -360
rect 1140 -372 1152 -360
rect 1164 -372 1176 -360
rect 1188 -372 1200 -360
rect 1212 -372 1224 -360
rect 1236 -372 1248 -360
rect 1260 -372 1272 -360
rect 1284 -372 1296 -360
rect 1308 -372 1320 -360
rect 1332 -372 1344 -360
rect 1356 -372 1368 -360
rect 1380 -372 1392 -360
rect 1404 -372 1416 -360
rect 1428 -372 1440 -360
rect 1452 -372 1464 -360
rect 1476 -372 1488 -360
rect 1500 -372 1512 -360
rect 1524 -372 1536 -360
rect 1548 -372 1560 -360
rect 1572 -372 1584 -360
rect 1596 -372 1608 -360
rect 1620 -372 1632 -360
rect 1644 -372 1656 -360
rect 1668 -372 1680 -360
rect 1692 -372 1704 -360
rect 1716 -372 1728 -360
rect 1740 -372 1752 -360
rect 1764 -372 1776 -360
rect 1788 -372 1800 -360
rect 1812 -372 1824 -360
rect 1836 -372 1848 -360
rect 1860 -372 1872 -360
rect 1884 -372 1896 -360
rect 1908 -372 1920 -360
rect 1932 -372 1944 -360
rect 1956 -372 1968 -360
rect 1980 -372 1992 -360
rect 2004 -372 2016 -360
rect 2028 -372 2040 -360
rect 2052 -372 2064 -360
rect 2076 -372 2088 -360
rect 2100 -372 2112 -360
rect 2124 -372 2136 -360
rect 2148 -372 2160 -360
rect 2172 -372 2184 -360
rect 2196 -372 2208 -360
rect 2220 -372 2232 -360
rect 2244 -372 2256 -360
rect 2268 -372 2280 -360
rect 2292 -372 2304 -360
rect 2316 -372 2328 -360
rect 2340 -372 2352 -360
rect 2364 -372 2376 -360
rect 2388 -372 2400 -360
rect 2412 -372 2424 -360
rect 2436 -372 2448 -360
rect 2460 -372 2472 -360
rect 2484 -372 2496 -360
rect 2508 -372 2520 -360
rect 2532 -372 2544 -360
rect 2556 -372 2568 -360
rect 2580 -372 2592 -360
rect 2604 -372 2616 -360
rect 2628 -372 2640 -360
rect 2652 -372 2664 -360
rect 2676 -372 2688 -360
rect 2700 -372 2712 -360
rect 2724 -372 2736 -360
rect 2748 -372 2760 -360
rect 2772 -372 2784 -360
rect 2796 -372 2808 -360
rect 2820 -372 2832 -360
rect 2844 -372 2856 -360
rect 2868 -372 2880 -360
rect 2892 -372 2904 -360
rect 2916 -372 2928 -360
rect 2940 -372 2952 -360
<< metal3 >>
rect -1044 588 -1032 648
rect -1044 534 -1032 552
rect -1044 516 -1032 528
rect -1044 384 -1032 396
rect -1104 346 -1032 348
rect -1104 320 -1102 346
rect -1094 320 -1054 346
rect -1046 320 -1032 346
rect -1104 318 -1032 320
rect -1104 310 -1032 312
rect -1104 302 -1078 310
rect -1070 302 -1032 310
rect -1104 300 -1032 302
rect -1104 292 -1032 294
rect -1104 266 -1102 292
rect -1094 266 -1054 292
rect -1046 266 -1032 292
rect -1104 264 -1032 266
rect -1044 216 -1032 228
rect -1044 168 -1032 180
rect -1044 120 -1032 132
rect -1044 72 -1032 84
rect -1104 34 -1032 36
rect -1104 8 -1102 34
rect -1094 8 -1054 34
rect -1046 8 -1032 34
rect -1104 6 -1032 8
rect -1104 -2 -1032 0
rect -1104 -10 -1078 -2
rect -1070 -10 -1032 -2
rect -1104 -12 -1032 -10
rect -1104 -20 -1032 -18
rect -1104 -46 -1102 -20
rect -1094 -46 -1054 -20
rect -1046 -46 -1032 -20
rect -1104 -48 -1032 -46
rect -1044 -168 -1032 -108
<< via3 >>
rect -1102 320 -1094 346
rect -1054 320 -1046 346
rect 168 324 180 348
rect 2016 324 2028 348
rect -1078 302 -1070 310
rect -744 300 -732 312
rect -672 300 -660 312
rect 336 300 348 312
rect 816 300 828 312
rect 888 300 900 312
rect 1296 300 1308 312
rect 1368 300 1380 312
rect 1848 300 1860 312
rect 2856 300 2868 312
rect 2928 300 2940 312
rect -1102 266 -1094 292
rect -1054 266 -1046 292
rect 168 264 180 288
rect 2016 264 2028 288
rect -792 216 -780 228
rect -624 216 -612 228
rect -432 216 -420 228
rect 576 216 588 228
rect 768 216 780 228
rect 936 216 948 228
rect 1248 216 1260 228
rect 1416 216 1428 228
rect 1608 216 1620 228
rect 2616 216 2628 228
rect 2808 216 2820 228
rect 2976 216 2988 228
rect -144 168 -132 180
rect -72 168 -60 180
rect 216 168 228 180
rect 288 168 300 180
rect 1896 168 1908 180
rect 1968 168 1980 180
rect 2256 168 2268 180
rect 2328 168 2340 180
rect -384 120 -372 132
rect -312 120 -300 132
rect 48 120 60 132
rect 96 120 108 132
rect 456 120 468 132
rect 528 120 540 132
rect 1656 120 1668 132
rect 1728 120 1740 132
rect 2088 120 2100 132
rect 2136 120 2148 132
rect 2496 120 2508 132
rect 2568 120 2580 132
rect -864 72 -852 84
rect -552 72 -540 84
rect -264 72 -252 84
rect 408 72 420 84
rect 696 72 708 84
rect 1008 72 1020 84
rect 1176 72 1188 84
rect 1488 72 1500 84
rect 1776 72 1788 84
rect 2448 72 2460 84
rect 2736 72 2748 84
rect 3048 72 3060 84
rect -1102 8 -1094 34
rect -1054 8 -1046 34
rect -24 12 -12 36
rect 2208 12 2220 36
rect -1078 -10 -1070 -2
rect -912 -12 -900 0
rect -504 -12 -492 0
rect -192 -12 -180 0
rect 648 -12 660 0
rect 1056 -12 1068 0
rect 1128 -12 1140 0
rect 1536 -12 1548 0
rect 2376 -12 2388 0
rect 2688 -12 2700 0
rect 3096 -12 3108 0
rect -1102 -46 -1094 -20
rect -1054 -46 -1046 -20
rect -24 -48 -12 -24
rect 2208 -48 2220 -24
<< metal4 >>
rect -1020 888 2988 900
rect -1104 744 -1092 756
rect -1104 696 -1092 732
rect -1104 346 -1092 684
rect -1104 320 -1102 346
rect -1094 320 -1092 346
rect -1104 292 -1092 320
rect -1104 266 -1102 292
rect -1094 266 -1092 292
rect -1104 264 -1092 266
rect -1080 720 -1068 756
rect -1080 310 -1068 708
rect -1080 302 -1078 310
rect -1070 302 -1068 310
rect -1080 264 -1068 302
rect -1056 744 -1044 756
rect -1056 696 -1044 732
rect -1020 744 -1008 888
rect 2976 744 2988 888
rect -1020 720 2988 744
rect -1020 708 -996 720
rect -984 708 -972 720
rect -960 708 -948 720
rect -936 708 -924 720
rect -912 708 -900 720
rect -888 708 -876 720
rect -864 708 -852 720
rect -840 708 -828 720
rect -816 708 -804 720
rect -792 708 -780 720
rect -768 708 -756 720
rect -744 708 -732 720
rect -720 708 -708 720
rect -696 708 -684 720
rect -672 708 -660 720
rect -648 708 -636 720
rect -624 708 -612 720
rect -600 708 -588 720
rect -576 708 -564 720
rect -552 708 -540 720
rect -528 708 -516 720
rect -504 708 -492 720
rect -480 708 -468 720
rect -456 708 -444 720
rect -432 708 -420 720
rect -408 708 -396 720
rect -384 708 -372 720
rect -360 708 -348 720
rect -336 708 -324 720
rect -312 708 -300 720
rect -288 708 -276 720
rect -264 708 -252 720
rect -240 708 -228 720
rect -216 708 -204 720
rect -192 708 -180 720
rect -168 708 -156 720
rect -144 708 -132 720
rect -120 708 -108 720
rect -96 708 -84 720
rect -72 708 -60 720
rect -48 708 -36 720
rect -24 708 -12 720
rect 0 708 12 720
rect 24 708 36 720
rect 48 708 60 720
rect 72 708 84 720
rect 96 708 108 720
rect 120 708 132 720
rect 144 708 156 720
rect 168 708 180 720
rect 192 708 204 720
rect 216 708 228 720
rect 240 708 252 720
rect 264 708 276 720
rect 288 708 300 720
rect 312 708 324 720
rect 336 708 348 720
rect 360 708 372 720
rect 384 708 396 720
rect 408 708 420 720
rect 432 708 444 720
rect 456 708 468 720
rect 480 708 492 720
rect 504 708 516 720
rect 528 708 540 720
rect 552 708 564 720
rect 576 708 588 720
rect 600 708 612 720
rect 624 708 636 720
rect 648 708 660 720
rect 672 708 684 720
rect 696 708 708 720
rect 720 708 732 720
rect 744 708 756 720
rect 768 708 780 720
rect 792 708 804 720
rect 816 708 828 720
rect 840 708 852 720
rect 864 708 876 720
rect 888 708 900 720
rect 912 708 924 720
rect 936 708 948 720
rect 960 708 972 720
rect 984 708 996 720
rect 1008 708 1020 720
rect 1032 708 1044 720
rect 1056 708 1068 720
rect 1080 708 1092 720
rect 1104 708 1116 720
rect 1128 708 1140 720
rect 1152 708 1164 720
rect 1176 708 1188 720
rect 1200 708 1212 720
rect 1224 708 1236 720
rect 1248 708 1260 720
rect 1272 708 1284 720
rect 1296 708 1308 720
rect 1320 708 1332 720
rect 1344 708 1356 720
rect 1368 708 1380 720
rect 1392 708 1404 720
rect 1416 708 1428 720
rect 1440 708 1452 720
rect 1464 708 1476 720
rect 1488 708 1500 720
rect 1512 708 1524 720
rect 1536 708 1548 720
rect 1560 708 1572 720
rect 1584 708 1596 720
rect 1608 708 1620 720
rect 1632 708 1644 720
rect 1656 708 1668 720
rect 1680 708 1692 720
rect 1704 708 1716 720
rect 1728 708 1740 720
rect 1752 708 1764 720
rect 1776 708 1788 720
rect 1800 708 1812 720
rect 1824 708 1836 720
rect 1848 708 1860 720
rect 1872 708 1884 720
rect 1896 708 1908 720
rect 1920 708 1932 720
rect 1944 708 1956 720
rect 1968 708 1980 720
rect 1992 708 2004 720
rect 2016 708 2028 720
rect 2040 708 2052 720
rect 2064 708 2076 720
rect 2088 708 2100 720
rect 2112 708 2124 720
rect 2136 708 2148 720
rect 2160 708 2172 720
rect 2184 708 2196 720
rect 2208 708 2220 720
rect 2232 708 2244 720
rect 2256 708 2268 720
rect 2280 708 2292 720
rect 2304 708 2316 720
rect 2328 708 2340 720
rect 2352 708 2364 720
rect 2376 708 2388 720
rect 2400 708 2412 720
rect 2424 708 2436 720
rect 2448 708 2460 720
rect 2472 708 2484 720
rect 2496 708 2508 720
rect 2520 708 2532 720
rect 2544 708 2556 720
rect 2568 708 2580 720
rect 2592 708 2604 720
rect 2616 708 2628 720
rect 2640 708 2652 720
rect 2664 708 2676 720
rect 2688 708 2700 720
rect 2712 708 2724 720
rect 2736 708 2748 720
rect 2760 708 2772 720
rect 2784 708 2796 720
rect 2808 708 2820 720
rect 2832 708 2844 720
rect 2856 708 2868 720
rect 2880 708 2892 720
rect 2904 708 2916 720
rect 2928 708 2940 720
rect 2952 708 2964 720
rect 2976 708 2988 720
rect -1020 684 2988 708
rect -1056 346 -1044 684
rect -1056 320 -1054 346
rect -1046 320 -1044 346
rect -1056 292 -1044 320
rect -1056 266 -1054 292
rect -1046 266 -1044 292
rect -1056 264 -1044 266
rect -1104 34 -1092 36
rect -1104 8 -1102 34
rect -1094 8 -1092 34
rect -1104 -20 -1092 8
rect -1104 -46 -1102 -20
rect -1094 -46 -1092 -20
rect -1104 -180 -1092 -46
rect -1104 -228 -1092 -192
rect -1104 -252 -1092 -240
rect -1080 -2 -1068 36
rect -1080 -10 -1078 -2
rect -1070 -10 -1068 -2
rect -1080 -204 -1068 -10
rect -1080 -252 -1068 -216
rect -1056 34 -1044 36
rect -1056 8 -1054 34
rect -1046 8 -1044 34
rect -1056 -20 -1044 8
rect -1056 -46 -1054 -20
rect -1046 -46 -1044 -20
rect -1056 -180 -1044 -46
rect -1056 -228 -1044 -192
rect -1056 -252 -1044 -240
rect -1020 -204 2988 -180
rect -1020 -216 -996 -204
rect -984 -216 -972 -204
rect -960 -216 -948 -204
rect -936 -216 -924 -204
rect -912 -216 -900 -204
rect -888 -216 -876 -204
rect -864 -216 -852 -204
rect -840 -216 -828 -204
rect -816 -216 -804 -204
rect -792 -216 -780 -204
rect -768 -216 -756 -204
rect -744 -216 -732 -204
rect -720 -216 -708 -204
rect -696 -216 -684 -204
rect -672 -216 -660 -204
rect -648 -216 -636 -204
rect -624 -216 -612 -204
rect -600 -216 -588 -204
rect -576 -216 -564 -204
rect -552 -216 -540 -204
rect -528 -216 -516 -204
rect -504 -216 -492 -204
rect -480 -216 -468 -204
rect -456 -216 -444 -204
rect -432 -216 -420 -204
rect -408 -216 -396 -204
rect -384 -216 -372 -204
rect -360 -216 -348 -204
rect -336 -216 -324 -204
rect -312 -216 -300 -204
rect -288 -216 -276 -204
rect -264 -216 -252 -204
rect -240 -216 -228 -204
rect -216 -216 -204 -204
rect -192 -216 -180 -204
rect -168 -216 -156 -204
rect -144 -216 -132 -204
rect -120 -216 -108 -204
rect -96 -216 -84 -204
rect -72 -216 -60 -204
rect -48 -216 -36 -204
rect -24 -216 -12 -204
rect 0 -216 12 -204
rect 24 -216 36 -204
rect 48 -216 60 -204
rect 72 -216 84 -204
rect 96 -216 108 -204
rect 120 -216 132 -204
rect 144 -216 156 -204
rect 168 -216 180 -204
rect 192 -216 204 -204
rect 216 -216 228 -204
rect 240 -216 252 -204
rect 264 -216 276 -204
rect 288 -216 300 -204
rect 312 -216 324 -204
rect 336 -216 348 -204
rect 360 -216 372 -204
rect 384 -216 396 -204
rect 408 -216 420 -204
rect 432 -216 444 -204
rect 456 -216 468 -204
rect 480 -216 492 -204
rect 504 -216 516 -204
rect 528 -216 540 -204
rect 552 -216 564 -204
rect 576 -216 588 -204
rect 600 -216 612 -204
rect 624 -216 636 -204
rect 648 -216 660 -204
rect 672 -216 684 -204
rect 696 -216 708 -204
rect 720 -216 732 -204
rect 744 -216 756 -204
rect 768 -216 780 -204
rect 792 -216 804 -204
rect 816 -216 828 -204
rect 840 -216 852 -204
rect 864 -216 876 -204
rect 888 -216 900 -204
rect 912 -216 924 -204
rect 936 -216 948 -204
rect 960 -216 972 -204
rect 984 -216 996 -204
rect 1008 -216 1020 -204
rect 1032 -216 1044 -204
rect 1056 -216 1068 -204
rect 1080 -216 1092 -204
rect 1104 -216 1116 -204
rect 1128 -216 1140 -204
rect 1152 -216 1164 -204
rect 1176 -216 1188 -204
rect 1200 -216 1212 -204
rect 1224 -216 1236 -204
rect 1248 -216 1260 -204
rect 1272 -216 1284 -204
rect 1296 -216 1308 -204
rect 1320 -216 1332 -204
rect 1344 -216 1356 -204
rect 1368 -216 1380 -204
rect 1392 -216 1404 -204
rect 1416 -216 1428 -204
rect 1440 -216 1452 -204
rect 1464 -216 1476 -204
rect 1488 -216 1500 -204
rect 1512 -216 1524 -204
rect 1536 -216 1548 -204
rect 1560 -216 1572 -204
rect 1584 -216 1596 -204
rect 1608 -216 1620 -204
rect 1632 -216 1644 -204
rect 1656 -216 1668 -204
rect 1680 -216 1692 -204
rect 1704 -216 1716 -204
rect 1728 -216 1740 -204
rect 1752 -216 1764 -204
rect 1776 -216 1788 -204
rect 1800 -216 1812 -204
rect 1824 -216 1836 -204
rect 1848 -216 1860 -204
rect 1872 -216 1884 -204
rect 1896 -216 1908 -204
rect 1920 -216 1932 -204
rect 1944 -216 1956 -204
rect 1968 -216 1980 -204
rect 1992 -216 2004 -204
rect 2016 -216 2028 -204
rect 2040 -216 2052 -204
rect 2064 -216 2076 -204
rect 2088 -216 2100 -204
rect 2112 -216 2124 -204
rect 2136 -216 2148 -204
rect 2160 -216 2172 -204
rect 2184 -216 2196 -204
rect 2208 -216 2220 -204
rect 2232 -216 2244 -204
rect 2256 -216 2268 -204
rect 2280 -216 2292 -204
rect 2304 -216 2316 -204
rect 2328 -216 2340 -204
rect 2352 -216 2364 -204
rect 2376 -216 2388 -204
rect 2400 -216 2412 -204
rect 2424 -216 2436 -204
rect 2448 -216 2460 -204
rect 2472 -216 2484 -204
rect 2496 -216 2508 -204
rect 2520 -216 2532 -204
rect 2544 -216 2556 -204
rect 2568 -216 2580 -204
rect 2592 -216 2604 -204
rect 2616 -216 2628 -204
rect 2640 -216 2652 -204
rect 2664 -216 2676 -204
rect 2688 -216 2700 -204
rect 2712 -216 2724 -204
rect 2736 -216 2748 -204
rect 2760 -216 2772 -204
rect 2784 -216 2796 -204
rect 2808 -216 2820 -204
rect 2832 -216 2844 -204
rect 2856 -216 2868 -204
rect 2880 -216 2892 -204
rect 2904 -216 2916 -204
rect 2928 -216 2940 -204
rect 2952 -216 2964 -204
rect 2976 -216 2988 -204
rect -1020 -240 2988 -216
rect -1020 -384 -1008 -240
rect 2976 -384 2988 -240
rect -1020 -396 2988 -384
<< via4 >>
rect -1104 732 -1092 744
rect -1104 684 -1092 696
rect -1080 708 -1068 720
rect -1056 732 -1044 744
rect -1056 684 -1044 696
rect -996 708 -984 720
rect -972 708 -960 720
rect -948 708 -936 720
rect -924 708 -912 720
rect -900 708 -888 720
rect -876 708 -864 720
rect -852 708 -840 720
rect -828 708 -816 720
rect -804 708 -792 720
rect -780 708 -768 720
rect -756 708 -744 720
rect -732 708 -720 720
rect -708 708 -696 720
rect -684 708 -672 720
rect -660 708 -648 720
rect -636 708 -624 720
rect -612 708 -600 720
rect -588 708 -576 720
rect -564 708 -552 720
rect -540 708 -528 720
rect -516 708 -504 720
rect -492 708 -480 720
rect -468 708 -456 720
rect -444 708 -432 720
rect -420 708 -408 720
rect -396 708 -384 720
rect -372 708 -360 720
rect -348 708 -336 720
rect -324 708 -312 720
rect -300 708 -288 720
rect -276 708 -264 720
rect -252 708 -240 720
rect -228 708 -216 720
rect -204 708 -192 720
rect -180 708 -168 720
rect -156 708 -144 720
rect -132 708 -120 720
rect -108 708 -96 720
rect -84 708 -72 720
rect -60 708 -48 720
rect -36 708 -24 720
rect -12 708 0 720
rect 12 708 24 720
rect 36 708 48 720
rect 60 708 72 720
rect 84 708 96 720
rect 108 708 120 720
rect 132 708 144 720
rect 156 708 168 720
rect 180 708 192 720
rect 204 708 216 720
rect 228 708 240 720
rect 252 708 264 720
rect 276 708 288 720
rect 300 708 312 720
rect 324 708 336 720
rect 348 708 360 720
rect 372 708 384 720
rect 396 708 408 720
rect 420 708 432 720
rect 444 708 456 720
rect 468 708 480 720
rect 492 708 504 720
rect 516 708 528 720
rect 540 708 552 720
rect 564 708 576 720
rect 588 708 600 720
rect 612 708 624 720
rect 636 708 648 720
rect 660 708 672 720
rect 684 708 696 720
rect 708 708 720 720
rect 732 708 744 720
rect 756 708 768 720
rect 780 708 792 720
rect 804 708 816 720
rect 828 708 840 720
rect 852 708 864 720
rect 876 708 888 720
rect 900 708 912 720
rect 924 708 936 720
rect 948 708 960 720
rect 972 708 984 720
rect 996 708 1008 720
rect 1020 708 1032 720
rect 1044 708 1056 720
rect 1068 708 1080 720
rect 1092 708 1104 720
rect 1116 708 1128 720
rect 1140 708 1152 720
rect 1164 708 1176 720
rect 1188 708 1200 720
rect 1212 708 1224 720
rect 1236 708 1248 720
rect 1260 708 1272 720
rect 1284 708 1296 720
rect 1308 708 1320 720
rect 1332 708 1344 720
rect 1356 708 1368 720
rect 1380 708 1392 720
rect 1404 708 1416 720
rect 1428 708 1440 720
rect 1452 708 1464 720
rect 1476 708 1488 720
rect 1500 708 1512 720
rect 1524 708 1536 720
rect 1548 708 1560 720
rect 1572 708 1584 720
rect 1596 708 1608 720
rect 1620 708 1632 720
rect 1644 708 1656 720
rect 1668 708 1680 720
rect 1692 708 1704 720
rect 1716 708 1728 720
rect 1740 708 1752 720
rect 1764 708 1776 720
rect 1788 708 1800 720
rect 1812 708 1824 720
rect 1836 708 1848 720
rect 1860 708 1872 720
rect 1884 708 1896 720
rect 1908 708 1920 720
rect 1932 708 1944 720
rect 1956 708 1968 720
rect 1980 708 1992 720
rect 2004 708 2016 720
rect 2028 708 2040 720
rect 2052 708 2064 720
rect 2076 708 2088 720
rect 2100 708 2112 720
rect 2124 708 2136 720
rect 2148 708 2160 720
rect 2172 708 2184 720
rect 2196 708 2208 720
rect 2220 708 2232 720
rect 2244 708 2256 720
rect 2268 708 2280 720
rect 2292 708 2304 720
rect 2316 708 2328 720
rect 2340 708 2352 720
rect 2364 708 2376 720
rect 2388 708 2400 720
rect 2412 708 2424 720
rect 2436 708 2448 720
rect 2460 708 2472 720
rect 2484 708 2496 720
rect 2508 708 2520 720
rect 2532 708 2544 720
rect 2556 708 2568 720
rect 2580 708 2592 720
rect 2604 708 2616 720
rect 2628 708 2640 720
rect 2652 708 2664 720
rect 2676 708 2688 720
rect 2700 708 2712 720
rect 2724 708 2736 720
rect 2748 708 2760 720
rect 2772 708 2784 720
rect 2796 708 2808 720
rect 2820 708 2832 720
rect 2844 708 2856 720
rect 2868 708 2880 720
rect 2892 708 2904 720
rect 2916 708 2928 720
rect 2940 708 2952 720
rect 2964 708 2976 720
rect -1104 -192 -1092 -180
rect -1104 -240 -1092 -228
rect -1080 -216 -1068 -204
rect -1056 -192 -1044 -180
rect -1056 -240 -1044 -228
rect -996 -216 -984 -204
rect -972 -216 -960 -204
rect -948 -216 -936 -204
rect -924 -216 -912 -204
rect -900 -216 -888 -204
rect -876 -216 -864 -204
rect -852 -216 -840 -204
rect -828 -216 -816 -204
rect -804 -216 -792 -204
rect -780 -216 -768 -204
rect -756 -216 -744 -204
rect -732 -216 -720 -204
rect -708 -216 -696 -204
rect -684 -216 -672 -204
rect -660 -216 -648 -204
rect -636 -216 -624 -204
rect -612 -216 -600 -204
rect -588 -216 -576 -204
rect -564 -216 -552 -204
rect -540 -216 -528 -204
rect -516 -216 -504 -204
rect -492 -216 -480 -204
rect -468 -216 -456 -204
rect -444 -216 -432 -204
rect -420 -216 -408 -204
rect -396 -216 -384 -204
rect -372 -216 -360 -204
rect -348 -216 -336 -204
rect -324 -216 -312 -204
rect -300 -216 -288 -204
rect -276 -216 -264 -204
rect -252 -216 -240 -204
rect -228 -216 -216 -204
rect -204 -216 -192 -204
rect -180 -216 -168 -204
rect -156 -216 -144 -204
rect -132 -216 -120 -204
rect -108 -216 -96 -204
rect -84 -216 -72 -204
rect -60 -216 -48 -204
rect -36 -216 -24 -204
rect -12 -216 0 -204
rect 12 -216 24 -204
rect 36 -216 48 -204
rect 60 -216 72 -204
rect 84 -216 96 -204
rect 108 -216 120 -204
rect 132 -216 144 -204
rect 156 -216 168 -204
rect 180 -216 192 -204
rect 204 -216 216 -204
rect 228 -216 240 -204
rect 252 -216 264 -204
rect 276 -216 288 -204
rect 300 -216 312 -204
rect 324 -216 336 -204
rect 348 -216 360 -204
rect 372 -216 384 -204
rect 396 -216 408 -204
rect 420 -216 432 -204
rect 444 -216 456 -204
rect 468 -216 480 -204
rect 492 -216 504 -204
rect 516 -216 528 -204
rect 540 -216 552 -204
rect 564 -216 576 -204
rect 588 -216 600 -204
rect 612 -216 624 -204
rect 636 -216 648 -204
rect 660 -216 672 -204
rect 684 -216 696 -204
rect 708 -216 720 -204
rect 732 -216 744 -204
rect 756 -216 768 -204
rect 780 -216 792 -204
rect 804 -216 816 -204
rect 828 -216 840 -204
rect 852 -216 864 -204
rect 876 -216 888 -204
rect 900 -216 912 -204
rect 924 -216 936 -204
rect 948 -216 960 -204
rect 972 -216 984 -204
rect 996 -216 1008 -204
rect 1020 -216 1032 -204
rect 1044 -216 1056 -204
rect 1068 -216 1080 -204
rect 1092 -216 1104 -204
rect 1116 -216 1128 -204
rect 1140 -216 1152 -204
rect 1164 -216 1176 -204
rect 1188 -216 1200 -204
rect 1212 -216 1224 -204
rect 1236 -216 1248 -204
rect 1260 -216 1272 -204
rect 1284 -216 1296 -204
rect 1308 -216 1320 -204
rect 1332 -216 1344 -204
rect 1356 -216 1368 -204
rect 1380 -216 1392 -204
rect 1404 -216 1416 -204
rect 1428 -216 1440 -204
rect 1452 -216 1464 -204
rect 1476 -216 1488 -204
rect 1500 -216 1512 -204
rect 1524 -216 1536 -204
rect 1548 -216 1560 -204
rect 1572 -216 1584 -204
rect 1596 -216 1608 -204
rect 1620 -216 1632 -204
rect 1644 -216 1656 -204
rect 1668 -216 1680 -204
rect 1692 -216 1704 -204
rect 1716 -216 1728 -204
rect 1740 -216 1752 -204
rect 1764 -216 1776 -204
rect 1788 -216 1800 -204
rect 1812 -216 1824 -204
rect 1836 -216 1848 -204
rect 1860 -216 1872 -204
rect 1884 -216 1896 -204
rect 1908 -216 1920 -204
rect 1932 -216 1944 -204
rect 1956 -216 1968 -204
rect 1980 -216 1992 -204
rect 2004 -216 2016 -204
rect 2028 -216 2040 -204
rect 2052 -216 2064 -204
rect 2076 -216 2088 -204
rect 2100 -216 2112 -204
rect 2124 -216 2136 -204
rect 2148 -216 2160 -204
rect 2172 -216 2184 -204
rect 2196 -216 2208 -204
rect 2220 -216 2232 -204
rect 2244 -216 2256 -204
rect 2268 -216 2280 -204
rect 2292 -216 2304 -204
rect 2316 -216 2328 -204
rect 2340 -216 2352 -204
rect 2364 -216 2376 -204
rect 2388 -216 2400 -204
rect 2412 -216 2424 -204
rect 2436 -216 2448 -204
rect 2460 -216 2472 -204
rect 2484 -216 2496 -204
rect 2508 -216 2520 -204
rect 2532 -216 2544 -204
rect 2556 -216 2568 -204
rect 2580 -216 2592 -204
rect 2604 -216 2616 -204
rect 2628 -216 2640 -204
rect 2652 -216 2664 -204
rect 2676 -216 2688 -204
rect 2700 -216 2712 -204
rect 2724 -216 2736 -204
rect 2748 -216 2760 -204
rect 2772 -216 2784 -204
rect 2796 -216 2808 -204
rect 2820 -216 2832 -204
rect 2844 -216 2856 -204
rect 2868 -216 2880 -204
rect 2892 -216 2904 -204
rect 2916 -216 2928 -204
rect 2940 -216 2952 -204
rect 2964 -216 2976 -204
<< metal5 >>
rect -1020 876 2988 900
rect -1020 864 -996 876
rect -984 864 -948 876
rect -936 864 -924 876
rect -912 864 -876 876
rect -864 864 -852 876
rect -840 864 -804 876
rect -792 864 -780 876
rect -768 864 -732 876
rect -720 864 -708 876
rect -696 864 -660 876
rect -648 864 -636 876
rect -624 864 -588 876
rect -576 864 -564 876
rect -552 864 -516 876
rect -504 864 -492 876
rect -480 864 -444 876
rect -432 864 -420 876
rect -408 864 -372 876
rect -360 864 -348 876
rect -336 864 -300 876
rect -288 864 -276 876
rect -264 864 -228 876
rect -216 864 -204 876
rect -192 864 -156 876
rect -144 864 -132 876
rect -120 864 -84 876
rect -72 864 -60 876
rect -48 864 -12 876
rect 0 864 12 876
rect 24 864 60 876
rect 72 864 84 876
rect 96 864 132 876
rect 144 864 156 876
rect 168 864 204 876
rect 216 864 228 876
rect 240 864 276 876
rect 288 864 300 876
rect 312 864 348 876
rect 360 864 372 876
rect 384 864 420 876
rect 432 864 444 876
rect 456 864 492 876
rect 504 864 516 876
rect 528 864 564 876
rect 576 864 588 876
rect 600 864 636 876
rect 648 864 660 876
rect 672 864 708 876
rect 720 864 732 876
rect 744 864 780 876
rect 792 864 804 876
rect 816 864 852 876
rect 864 864 876 876
rect 888 864 924 876
rect 936 864 948 876
rect 960 864 996 876
rect 1008 864 1020 876
rect 1032 864 1068 876
rect 1080 864 1092 876
rect 1104 864 1140 876
rect 1152 864 1164 876
rect 1176 864 1212 876
rect 1224 864 1236 876
rect 1248 864 1284 876
rect 1296 864 1308 876
rect 1320 864 1356 876
rect 1368 864 1380 876
rect 1392 864 1428 876
rect 1440 864 1452 876
rect 1464 864 1500 876
rect 1512 864 1524 876
rect 1536 864 1572 876
rect 1584 864 1596 876
rect 1608 864 1644 876
rect 1656 864 1668 876
rect 1680 864 1716 876
rect 1728 864 1740 876
rect 1752 864 1788 876
rect 1800 864 1812 876
rect 1824 864 1860 876
rect 1872 864 1884 876
rect 1896 864 1932 876
rect 1944 864 1956 876
rect 1968 864 2004 876
rect 2016 864 2028 876
rect 2040 864 2076 876
rect 2088 864 2100 876
rect 2112 864 2148 876
rect 2160 864 2172 876
rect 2184 864 2220 876
rect 2232 864 2244 876
rect 2256 864 2292 876
rect 2304 864 2316 876
rect 2328 864 2364 876
rect 2376 864 2388 876
rect 2400 864 2436 876
rect 2448 864 2460 876
rect 2472 864 2484 876
rect 2496 864 2532 876
rect 2544 864 2556 876
rect 2568 864 2604 876
rect 2616 864 2628 876
rect 2640 864 2676 876
rect 2688 864 2700 876
rect 2712 864 2724 876
rect 2736 864 2772 876
rect 2784 864 2796 876
rect 2808 864 2844 876
rect 2856 864 2868 876
rect 2880 864 2916 876
rect 2928 864 2940 876
rect 2952 864 2988 876
rect -1020 840 2988 864
rect -1020 828 -996 840
rect -984 828 -972 840
rect -960 828 -948 840
rect -936 828 -924 840
rect -912 828 -900 840
rect -888 828 -876 840
rect -864 828 -852 840
rect -840 828 -828 840
rect -816 828 -804 840
rect -792 828 -780 840
rect -768 828 -756 840
rect -744 828 -732 840
rect -720 828 -708 840
rect -696 828 -684 840
rect -672 828 -660 840
rect -648 828 -636 840
rect -624 828 -612 840
rect -600 828 -588 840
rect -576 828 -564 840
rect -552 828 -540 840
rect -528 828 -516 840
rect -504 828 -492 840
rect -480 828 -468 840
rect -456 828 -444 840
rect -432 828 -420 840
rect -408 828 -396 840
rect -384 828 -372 840
rect -360 828 -348 840
rect -336 828 -324 840
rect -312 828 -300 840
rect -288 828 -276 840
rect -264 828 -252 840
rect -240 828 -228 840
rect -216 828 -204 840
rect -192 828 -180 840
rect -168 828 -156 840
rect -144 828 -132 840
rect -120 828 -108 840
rect -96 828 -84 840
rect -72 828 -60 840
rect -48 828 -36 840
rect -24 828 -12 840
rect 0 828 12 840
rect 24 828 36 840
rect 48 828 60 840
rect 72 828 84 840
rect 96 828 108 840
rect 120 828 132 840
rect 144 828 156 840
rect 168 828 180 840
rect 192 828 204 840
rect 216 828 228 840
rect 240 828 252 840
rect 264 828 276 840
rect 288 828 300 840
rect 312 828 324 840
rect 336 828 348 840
rect 360 828 372 840
rect 384 828 396 840
rect 408 828 420 840
rect 432 828 444 840
rect 456 828 468 840
rect 480 828 492 840
rect 504 828 516 840
rect 528 828 540 840
rect 552 828 564 840
rect 576 828 588 840
rect 600 828 612 840
rect 624 828 636 840
rect 648 828 660 840
rect 672 828 684 840
rect 696 828 708 840
rect 720 828 732 840
rect 744 828 756 840
rect 768 828 780 840
rect 792 828 804 840
rect 816 828 828 840
rect 840 828 852 840
rect 864 828 876 840
rect 888 828 900 840
rect 912 828 924 840
rect 936 828 948 840
rect 960 828 972 840
rect 984 828 996 840
rect 1008 828 1020 840
rect 1032 828 1044 840
rect 1056 828 1068 840
rect 1080 828 1092 840
rect 1104 828 1116 840
rect 1128 828 1140 840
rect 1152 828 1164 840
rect 1176 828 1188 840
rect 1200 828 1212 840
rect 1224 828 1236 840
rect 1248 828 1260 840
rect 1272 828 1284 840
rect 1296 828 1308 840
rect 1320 828 1332 840
rect 1344 828 1356 840
rect 1368 828 1380 840
rect 1392 828 1404 840
rect 1416 828 1428 840
rect 1440 828 1452 840
rect 1464 828 1476 840
rect 1488 828 1500 840
rect 1512 828 1524 840
rect 1536 828 1548 840
rect 1560 828 1572 840
rect 1584 828 1596 840
rect 1608 828 1620 840
rect 1632 828 1644 840
rect 1656 828 1668 840
rect 1680 828 1692 840
rect 1704 828 1716 840
rect 1728 828 1740 840
rect 1752 828 1764 840
rect 1776 828 1788 840
rect 1800 828 1812 840
rect 1824 828 1836 840
rect 1848 828 1860 840
rect 1872 828 1884 840
rect 1896 828 1908 840
rect 1920 828 1932 840
rect 1944 828 1956 840
rect 1968 828 1980 840
rect 1992 828 2004 840
rect 2016 828 2028 840
rect 2040 828 2052 840
rect 2064 828 2076 840
rect 2088 828 2100 840
rect 2112 828 2124 840
rect 2136 828 2148 840
rect 2160 828 2172 840
rect 2184 828 2196 840
rect 2208 828 2220 840
rect 2232 828 2244 840
rect 2256 828 2268 840
rect 2280 828 2292 840
rect 2304 828 2316 840
rect 2328 828 2340 840
rect 2352 828 2364 840
rect 2376 828 2388 840
rect 2400 828 2412 840
rect 2424 828 2436 840
rect 2448 828 2460 840
rect 2472 828 2484 840
rect 2496 828 2508 840
rect 2520 828 2532 840
rect 2544 828 2556 840
rect 2568 828 2580 840
rect 2592 828 2604 840
rect 2616 828 2628 840
rect 2640 828 2652 840
rect 2664 828 2676 840
rect 2688 828 2700 840
rect 2712 828 2724 840
rect 2736 828 2748 840
rect 2760 828 2772 840
rect 2784 828 2796 840
rect 2808 828 2820 840
rect 2832 828 2844 840
rect 2856 828 2868 840
rect 2880 828 2892 840
rect 2904 828 2916 840
rect 2928 828 2940 840
rect 2952 828 2988 840
rect -1020 804 2988 828
rect -1020 792 -996 804
rect -984 792 -972 804
rect -960 792 -948 804
rect -936 792 -924 804
rect -912 792 -900 804
rect -888 792 -876 804
rect -864 792 -852 804
rect -840 792 -828 804
rect -816 792 -804 804
rect -792 792 -780 804
rect -768 792 -756 804
rect -744 792 -732 804
rect -720 792 -708 804
rect -696 792 -684 804
rect -672 792 -660 804
rect -648 792 -636 804
rect -624 792 -612 804
rect -600 792 -588 804
rect -576 792 -564 804
rect -552 792 -540 804
rect -528 792 -516 804
rect -504 792 -492 804
rect -480 792 -468 804
rect -456 792 -444 804
rect -432 792 -420 804
rect -408 792 -396 804
rect -384 792 -372 804
rect -360 792 -348 804
rect -336 792 -324 804
rect -312 792 -300 804
rect -288 792 -276 804
rect -264 792 -252 804
rect -240 792 -228 804
rect -216 792 -204 804
rect -192 792 -180 804
rect -168 792 -156 804
rect -144 792 -132 804
rect -120 792 -108 804
rect -96 792 -84 804
rect -72 792 -60 804
rect -48 792 -36 804
rect -24 792 -12 804
rect 0 792 12 804
rect 24 792 36 804
rect 48 792 60 804
rect 72 792 84 804
rect 96 792 108 804
rect 120 792 132 804
rect 144 792 156 804
rect 168 792 180 804
rect 192 792 204 804
rect 216 792 228 804
rect 240 792 252 804
rect 264 792 276 804
rect 288 792 300 804
rect 312 792 324 804
rect 336 792 348 804
rect 360 792 372 804
rect 384 792 396 804
rect 408 792 420 804
rect 432 792 444 804
rect 456 792 468 804
rect 480 792 492 804
rect 504 792 516 804
rect 528 792 540 804
rect 552 792 564 804
rect 576 792 588 804
rect 600 792 612 804
rect 624 792 636 804
rect 648 792 660 804
rect 672 792 684 804
rect 696 792 708 804
rect 720 792 732 804
rect 744 792 756 804
rect 768 792 780 804
rect 792 792 804 804
rect 816 792 828 804
rect 840 792 852 804
rect 864 792 876 804
rect 888 792 900 804
rect 912 792 924 804
rect 936 792 948 804
rect 960 792 972 804
rect 984 792 996 804
rect 1008 792 1020 804
rect 1032 792 1044 804
rect 1056 792 1068 804
rect 1080 792 1092 804
rect 1104 792 1116 804
rect 1128 792 1140 804
rect 1152 792 1164 804
rect 1176 792 1188 804
rect 1200 792 1212 804
rect 1224 792 1236 804
rect 1248 792 1260 804
rect 1272 792 1284 804
rect 1296 792 1308 804
rect 1320 792 1332 804
rect 1344 792 1356 804
rect 1368 792 1380 804
rect 1392 792 1404 804
rect 1416 792 1428 804
rect 1440 792 1452 804
rect 1464 792 1476 804
rect 1488 792 1500 804
rect 1512 792 1524 804
rect 1536 792 1548 804
rect 1560 792 1572 804
rect 1584 792 1596 804
rect 1608 792 1620 804
rect 1632 792 1644 804
rect 1656 792 1668 804
rect 1680 792 1692 804
rect 1704 792 1716 804
rect 1728 792 1740 804
rect 1752 792 1764 804
rect 1776 792 1788 804
rect 1800 792 1812 804
rect 1824 792 1836 804
rect 1848 792 1860 804
rect 1872 792 1884 804
rect 1896 792 1908 804
rect 1920 792 1932 804
rect 1944 792 1956 804
rect 1968 792 1980 804
rect 1992 792 2004 804
rect 2016 792 2028 804
rect 2040 792 2052 804
rect 2064 792 2076 804
rect 2088 792 2100 804
rect 2112 792 2124 804
rect 2136 792 2148 804
rect 2160 792 2172 804
rect 2184 792 2196 804
rect 2208 792 2220 804
rect 2232 792 2244 804
rect 2256 792 2268 804
rect 2280 792 2292 804
rect 2304 792 2316 804
rect 2328 792 2340 804
rect 2352 792 2364 804
rect 2376 792 2388 804
rect 2400 792 2412 804
rect 2424 792 2436 804
rect 2448 792 2460 804
rect 2472 792 2484 804
rect 2496 792 2508 804
rect 2520 792 2532 804
rect 2544 792 2556 804
rect 2568 792 2580 804
rect 2592 792 2604 804
rect 2616 792 2628 804
rect 2640 792 2652 804
rect 2664 792 2676 804
rect 2688 792 2700 804
rect 2712 792 2724 804
rect 2736 792 2748 804
rect 2760 792 2772 804
rect 2784 792 2796 804
rect 2808 792 2820 804
rect 2832 792 2844 804
rect 2856 792 2868 804
rect 2880 792 2892 804
rect 2904 792 2916 804
rect 2928 792 2940 804
rect 2952 792 2988 804
rect -1020 768 2988 792
rect -1020 756 -996 768
rect -984 756 -972 768
rect -960 756 -948 768
rect -936 756 -924 768
rect -912 756 -900 768
rect -888 756 -876 768
rect -864 756 -852 768
rect -840 756 -828 768
rect -816 756 -804 768
rect -792 756 -780 768
rect -768 756 -756 768
rect -744 756 -732 768
rect -720 756 -708 768
rect -696 756 -684 768
rect -672 756 -660 768
rect -648 756 -636 768
rect -624 756 -612 768
rect -600 756 -588 768
rect -576 756 -564 768
rect -552 756 -540 768
rect -528 756 -516 768
rect -504 756 -492 768
rect -480 756 -468 768
rect -456 756 -444 768
rect -432 756 -420 768
rect -408 756 -396 768
rect -384 756 -372 768
rect -360 756 -348 768
rect -336 756 -324 768
rect -312 756 -300 768
rect -288 756 -276 768
rect -264 756 -252 768
rect -240 756 -228 768
rect -216 756 -204 768
rect -192 756 -180 768
rect -168 756 -156 768
rect -144 756 -132 768
rect -120 756 -108 768
rect -96 756 -84 768
rect -72 756 -60 768
rect -48 756 -36 768
rect -24 756 -12 768
rect 0 756 12 768
rect 24 756 36 768
rect 48 756 60 768
rect 72 756 84 768
rect 96 756 108 768
rect 120 756 132 768
rect 144 756 156 768
rect 168 756 180 768
rect 192 756 204 768
rect 216 756 228 768
rect 240 756 252 768
rect 264 756 276 768
rect 288 756 300 768
rect 312 756 324 768
rect 336 756 348 768
rect 360 756 372 768
rect 384 756 396 768
rect 408 756 420 768
rect 432 756 444 768
rect 456 756 468 768
rect 480 756 492 768
rect 504 756 516 768
rect 528 756 540 768
rect 552 756 564 768
rect 576 756 588 768
rect 600 756 612 768
rect 624 756 636 768
rect 648 756 660 768
rect 672 756 684 768
rect 696 756 708 768
rect 720 756 732 768
rect 744 756 756 768
rect 768 756 780 768
rect 792 756 804 768
rect 816 756 828 768
rect 840 756 852 768
rect 864 756 876 768
rect 888 756 900 768
rect 912 756 924 768
rect 936 756 948 768
rect 960 756 972 768
rect 984 756 996 768
rect 1008 756 1020 768
rect 1032 756 1044 768
rect 1056 756 1068 768
rect 1080 756 1092 768
rect 1104 756 1116 768
rect 1128 756 1140 768
rect 1152 756 1164 768
rect 1176 756 1188 768
rect 1200 756 1212 768
rect 1224 756 1236 768
rect 1248 756 1260 768
rect 1272 756 1284 768
rect 1296 756 1308 768
rect 1320 756 1332 768
rect 1344 756 1356 768
rect 1368 756 1380 768
rect 1392 756 1404 768
rect 1416 756 1428 768
rect 1440 756 1452 768
rect 1464 756 1476 768
rect 1488 756 1500 768
rect 1512 756 1524 768
rect 1536 756 1548 768
rect 1560 756 1572 768
rect 1584 756 1596 768
rect 1608 756 1620 768
rect 1632 756 1644 768
rect 1656 756 1668 768
rect 1680 756 1692 768
rect 1704 756 1716 768
rect 1728 756 1740 768
rect 1752 756 1764 768
rect 1776 756 1788 768
rect 1800 756 1812 768
rect 1824 756 1836 768
rect 1848 756 1860 768
rect 1872 756 1884 768
rect 1896 756 1908 768
rect 1920 756 1932 768
rect 1944 756 1956 768
rect 1968 756 1980 768
rect 1992 756 2004 768
rect 2016 756 2028 768
rect 2040 756 2052 768
rect 2064 756 2076 768
rect 2088 756 2100 768
rect 2112 756 2124 768
rect 2136 756 2148 768
rect 2160 756 2172 768
rect 2184 756 2196 768
rect 2208 756 2220 768
rect 2232 756 2244 768
rect 2256 756 2268 768
rect 2280 756 2292 768
rect 2304 756 2316 768
rect 2328 756 2340 768
rect 2352 756 2364 768
rect 2376 756 2388 768
rect 2400 756 2412 768
rect 2424 756 2436 768
rect 2448 756 2460 768
rect 2472 756 2484 768
rect 2496 756 2508 768
rect 2520 756 2532 768
rect 2544 756 2556 768
rect 2568 756 2580 768
rect 2592 756 2604 768
rect 2616 756 2628 768
rect 2640 756 2652 768
rect 2664 756 2676 768
rect 2688 756 2700 768
rect 2712 756 2724 768
rect 2736 756 2748 768
rect 2760 756 2772 768
rect 2784 756 2796 768
rect 2808 756 2820 768
rect 2832 756 2844 768
rect 2856 756 2868 768
rect 2880 756 2892 768
rect 2904 756 2916 768
rect 2928 756 2940 768
rect 2952 756 2988 768
rect -1020 744 2988 756
rect -1116 732 -1104 744
rect -1092 732 -1056 744
rect -1044 732 2988 744
rect -1116 708 -1080 720
rect -1068 708 -996 720
rect -984 708 -972 720
rect -960 708 -948 720
rect -936 708 -924 720
rect -912 708 -900 720
rect -888 708 -876 720
rect -864 708 -852 720
rect -840 708 -828 720
rect -816 708 -804 720
rect -792 708 -780 720
rect -768 708 -756 720
rect -744 708 -732 720
rect -720 708 -708 720
rect -696 708 -684 720
rect -672 708 -660 720
rect -648 708 -636 720
rect -624 708 -612 720
rect -600 708 -588 720
rect -576 708 -564 720
rect -552 708 -540 720
rect -528 708 -516 720
rect -504 708 -492 720
rect -480 708 -468 720
rect -456 708 -444 720
rect -432 708 -420 720
rect -408 708 -396 720
rect -384 708 -372 720
rect -360 708 -348 720
rect -336 708 -324 720
rect -312 708 -300 720
rect -288 708 -276 720
rect -264 708 -252 720
rect -240 708 -228 720
rect -216 708 -204 720
rect -192 708 -180 720
rect -168 708 -156 720
rect -144 708 -132 720
rect -120 708 -108 720
rect -96 708 -84 720
rect -72 708 -60 720
rect -48 708 -36 720
rect -24 708 -12 720
rect 0 708 12 720
rect 24 708 36 720
rect 48 708 60 720
rect 72 708 84 720
rect 96 708 108 720
rect 120 708 132 720
rect 144 708 156 720
rect 168 708 180 720
rect 192 708 204 720
rect 216 708 228 720
rect 240 708 252 720
rect 264 708 276 720
rect 288 708 300 720
rect 312 708 324 720
rect 336 708 348 720
rect 360 708 372 720
rect 384 708 396 720
rect 408 708 420 720
rect 432 708 444 720
rect 456 708 468 720
rect 480 708 492 720
rect 504 708 516 720
rect 528 708 540 720
rect 552 708 564 720
rect 576 708 588 720
rect 600 708 612 720
rect 624 708 636 720
rect 648 708 660 720
rect 672 708 684 720
rect 696 708 708 720
rect 720 708 732 720
rect 744 708 756 720
rect 768 708 780 720
rect 792 708 804 720
rect 816 708 828 720
rect 840 708 852 720
rect 864 708 876 720
rect 888 708 900 720
rect 912 708 924 720
rect 936 708 948 720
rect 960 708 972 720
rect 984 708 996 720
rect 1008 708 1020 720
rect 1032 708 1044 720
rect 1056 708 1068 720
rect 1080 708 1092 720
rect 1104 708 1116 720
rect 1128 708 1140 720
rect 1152 708 1164 720
rect 1176 708 1188 720
rect 1200 708 1212 720
rect 1224 708 1236 720
rect 1248 708 1260 720
rect 1272 708 1284 720
rect 1296 708 1308 720
rect 1320 708 1332 720
rect 1344 708 1356 720
rect 1368 708 1380 720
rect 1392 708 1404 720
rect 1416 708 1428 720
rect 1440 708 1452 720
rect 1464 708 1476 720
rect 1488 708 1500 720
rect 1512 708 1524 720
rect 1536 708 1548 720
rect 1560 708 1572 720
rect 1584 708 1596 720
rect 1608 708 1620 720
rect 1632 708 1644 720
rect 1656 708 1668 720
rect 1680 708 1692 720
rect 1704 708 1716 720
rect 1728 708 1740 720
rect 1752 708 1764 720
rect 1776 708 1788 720
rect 1800 708 1812 720
rect 1824 708 1836 720
rect 1848 708 1860 720
rect 1872 708 1884 720
rect 1896 708 1908 720
rect 1920 708 1932 720
rect 1944 708 1956 720
rect 1968 708 1980 720
rect 1992 708 2004 720
rect 2016 708 2028 720
rect 2040 708 2052 720
rect 2064 708 2076 720
rect 2088 708 2100 720
rect 2112 708 2124 720
rect 2136 708 2148 720
rect 2160 708 2172 720
rect 2184 708 2196 720
rect 2208 708 2220 720
rect 2232 708 2244 720
rect 2256 708 2268 720
rect 2280 708 2292 720
rect 2304 708 2316 720
rect 2328 708 2340 720
rect 2352 708 2364 720
rect 2376 708 2388 720
rect 2400 708 2412 720
rect 2424 708 2436 720
rect 2448 708 2460 720
rect 2472 708 2484 720
rect 2496 708 2508 720
rect 2520 708 2532 720
rect 2544 708 2556 720
rect 2568 708 2580 720
rect 2592 708 2604 720
rect 2616 708 2628 720
rect 2640 708 2652 720
rect 2664 708 2676 720
rect 2688 708 2700 720
rect 2712 708 2724 720
rect 2736 708 2748 720
rect 2760 708 2772 720
rect 2784 708 2796 720
rect 2808 708 2820 720
rect 2832 708 2844 720
rect 2856 708 2868 720
rect 2880 708 2892 720
rect 2904 708 2916 720
rect 2928 708 2940 720
rect 2952 708 2964 720
rect 2976 708 2988 720
rect -1116 684 -1104 696
rect -1092 684 -1056 696
rect -1044 684 2988 696
rect -1116 -192 -1104 -180
rect -1092 -192 -1056 -180
rect -1044 -192 2988 -180
rect -1116 -216 -1080 -204
rect -1068 -216 -996 -204
rect -984 -216 -972 -204
rect -960 -216 -948 -204
rect -936 -216 -924 -204
rect -912 -216 -900 -204
rect -888 -216 -876 -204
rect -864 -216 -852 -204
rect -840 -216 -828 -204
rect -816 -216 -804 -204
rect -792 -216 -780 -204
rect -768 -216 -756 -204
rect -744 -216 -732 -204
rect -720 -216 -708 -204
rect -696 -216 -684 -204
rect -672 -216 -660 -204
rect -648 -216 -636 -204
rect -624 -216 -612 -204
rect -600 -216 -588 -204
rect -576 -216 -564 -204
rect -552 -216 -540 -204
rect -528 -216 -516 -204
rect -504 -216 -492 -204
rect -480 -216 -468 -204
rect -456 -216 -444 -204
rect -432 -216 -420 -204
rect -408 -216 -396 -204
rect -384 -216 -372 -204
rect -360 -216 -348 -204
rect -336 -216 -324 -204
rect -312 -216 -300 -204
rect -288 -216 -276 -204
rect -264 -216 -252 -204
rect -240 -216 -228 -204
rect -216 -216 -204 -204
rect -192 -216 -180 -204
rect -168 -216 -156 -204
rect -144 -216 -132 -204
rect -120 -216 -108 -204
rect -96 -216 -84 -204
rect -72 -216 -60 -204
rect -48 -216 -36 -204
rect -24 -216 -12 -204
rect 0 -216 12 -204
rect 24 -216 36 -204
rect 48 -216 60 -204
rect 72 -216 84 -204
rect 96 -216 108 -204
rect 120 -216 132 -204
rect 144 -216 156 -204
rect 168 -216 180 -204
rect 192 -216 204 -204
rect 216 -216 228 -204
rect 240 -216 252 -204
rect 264 -216 276 -204
rect 288 -216 300 -204
rect 312 -216 324 -204
rect 336 -216 348 -204
rect 360 -216 372 -204
rect 384 -216 396 -204
rect 408 -216 420 -204
rect 432 -216 444 -204
rect 456 -216 468 -204
rect 480 -216 492 -204
rect 504 -216 516 -204
rect 528 -216 540 -204
rect 552 -216 564 -204
rect 576 -216 588 -204
rect 600 -216 612 -204
rect 624 -216 636 -204
rect 648 -216 660 -204
rect 672 -216 684 -204
rect 696 -216 708 -204
rect 720 -216 732 -204
rect 744 -216 756 -204
rect 768 -216 780 -204
rect 792 -216 804 -204
rect 816 -216 828 -204
rect 840 -216 852 -204
rect 864 -216 876 -204
rect 888 -216 900 -204
rect 912 -216 924 -204
rect 936 -216 948 -204
rect 960 -216 972 -204
rect 984 -216 996 -204
rect 1008 -216 1020 -204
rect 1032 -216 1044 -204
rect 1056 -216 1068 -204
rect 1080 -216 1092 -204
rect 1104 -216 1116 -204
rect 1128 -216 1140 -204
rect 1152 -216 1164 -204
rect 1176 -216 1188 -204
rect 1200 -216 1212 -204
rect 1224 -216 1236 -204
rect 1248 -216 1260 -204
rect 1272 -216 1284 -204
rect 1296 -216 1308 -204
rect 1320 -216 1332 -204
rect 1344 -216 1356 -204
rect 1368 -216 1380 -204
rect 1392 -216 1404 -204
rect 1416 -216 1428 -204
rect 1440 -216 1452 -204
rect 1464 -216 1476 -204
rect 1488 -216 1500 -204
rect 1512 -216 1524 -204
rect 1536 -216 1548 -204
rect 1560 -216 1572 -204
rect 1584 -216 1596 -204
rect 1608 -216 1620 -204
rect 1632 -216 1644 -204
rect 1656 -216 1668 -204
rect 1680 -216 1692 -204
rect 1704 -216 1716 -204
rect 1728 -216 1740 -204
rect 1752 -216 1764 -204
rect 1776 -216 1788 -204
rect 1800 -216 1812 -204
rect 1824 -216 1836 -204
rect 1848 -216 1860 -204
rect 1872 -216 1884 -204
rect 1896 -216 1908 -204
rect 1920 -216 1932 -204
rect 1944 -216 1956 -204
rect 1968 -216 1980 -204
rect 1992 -216 2004 -204
rect 2016 -216 2028 -204
rect 2040 -216 2052 -204
rect 2064 -216 2076 -204
rect 2088 -216 2100 -204
rect 2112 -216 2124 -204
rect 2136 -216 2148 -204
rect 2160 -216 2172 -204
rect 2184 -216 2196 -204
rect 2208 -216 2220 -204
rect 2232 -216 2244 -204
rect 2256 -216 2268 -204
rect 2280 -216 2292 -204
rect 2304 -216 2316 -204
rect 2328 -216 2340 -204
rect 2352 -216 2364 -204
rect 2376 -216 2388 -204
rect 2400 -216 2412 -204
rect 2424 -216 2436 -204
rect 2448 -216 2460 -204
rect 2472 -216 2484 -204
rect 2496 -216 2508 -204
rect 2520 -216 2532 -204
rect 2544 -216 2556 -204
rect 2568 -216 2580 -204
rect 2592 -216 2604 -204
rect 2616 -216 2628 -204
rect 2640 -216 2652 -204
rect 2664 -216 2676 -204
rect 2688 -216 2700 -204
rect 2712 -216 2724 -204
rect 2736 -216 2748 -204
rect 2760 -216 2772 -204
rect 2784 -216 2796 -204
rect 2808 -216 2820 -204
rect 2832 -216 2844 -204
rect 2856 -216 2868 -204
rect 2880 -216 2892 -204
rect 2904 -216 2916 -204
rect 2928 -216 2940 -204
rect 2952 -216 2964 -204
rect 2976 -216 2988 -204
rect -1116 -240 -1104 -228
rect -1092 -240 -1056 -228
rect -1044 -240 2988 -228
rect -1020 -252 2988 -240
rect -1020 -264 -996 -252
rect -984 -264 -948 -252
rect -936 -264 -924 -252
rect -912 -264 -876 -252
rect -864 -264 -852 -252
rect -840 -264 -804 -252
rect -792 -264 -780 -252
rect -768 -264 -732 -252
rect -720 -264 -708 -252
rect -696 -264 -660 -252
rect -648 -264 -636 -252
rect -624 -264 -588 -252
rect -576 -264 -564 -252
rect -552 -264 -516 -252
rect -504 -264 -492 -252
rect -480 -264 -444 -252
rect -432 -264 -420 -252
rect -408 -264 -372 -252
rect -360 -264 -348 -252
rect -336 -264 -300 -252
rect -288 -264 -276 -252
rect -264 -264 -228 -252
rect -216 -264 -204 -252
rect -192 -264 -156 -252
rect -144 -264 -132 -252
rect -120 -264 -84 -252
rect -72 -264 -60 -252
rect -48 -264 -12 -252
rect 0 -264 12 -252
rect 24 -264 60 -252
rect 72 -264 84 -252
rect 96 -264 132 -252
rect 144 -264 156 -252
rect 168 -264 204 -252
rect 216 -264 228 -252
rect 240 -264 276 -252
rect 288 -264 300 -252
rect 312 -264 348 -252
rect 360 -264 372 -252
rect 384 -264 420 -252
rect 432 -264 444 -252
rect 456 -264 492 -252
rect 504 -264 516 -252
rect 528 -264 564 -252
rect 576 -264 588 -252
rect 600 -264 636 -252
rect 648 -264 660 -252
rect 672 -264 708 -252
rect 720 -264 732 -252
rect 744 -264 780 -252
rect 792 -264 804 -252
rect 816 -264 852 -252
rect 864 -264 876 -252
rect 888 -264 924 -252
rect 936 -264 948 -252
rect 960 -264 996 -252
rect 1008 -264 1020 -252
rect 1032 -264 1068 -252
rect 1080 -264 1092 -252
rect 1104 -264 1140 -252
rect 1152 -264 1164 -252
rect 1176 -264 1212 -252
rect 1224 -264 1236 -252
rect 1248 -264 1284 -252
rect 1296 -264 1308 -252
rect 1320 -264 1356 -252
rect 1368 -264 1380 -252
rect 1392 -264 1428 -252
rect 1440 -264 1452 -252
rect 1464 -264 1500 -252
rect 1512 -264 1524 -252
rect 1536 -264 1572 -252
rect 1584 -264 1596 -252
rect 1608 -264 1644 -252
rect 1656 -264 1668 -252
rect 1680 -264 1716 -252
rect 1728 -264 1740 -252
rect 1752 -264 1788 -252
rect 1800 -264 1812 -252
rect 1824 -264 1860 -252
rect 1872 -264 1884 -252
rect 1896 -264 1932 -252
rect 1944 -264 1956 -252
rect 1968 -264 2004 -252
rect 2016 -264 2028 -252
rect 2040 -264 2076 -252
rect 2088 -264 2100 -252
rect 2112 -264 2148 -252
rect 2160 -264 2172 -252
rect 2184 -264 2220 -252
rect 2232 -264 2244 -252
rect 2256 -264 2292 -252
rect 2304 -264 2316 -252
rect 2328 -264 2364 -252
rect 2376 -264 2388 -252
rect 2400 -264 2436 -252
rect 2448 -264 2460 -252
rect 2472 -264 2484 -252
rect 2496 -264 2532 -252
rect 2544 -264 2556 -252
rect 2568 -264 2604 -252
rect 2616 -264 2628 -252
rect 2640 -264 2676 -252
rect 2688 -264 2700 -252
rect 2712 -264 2724 -252
rect 2736 -264 2772 -252
rect 2784 -264 2796 -252
rect 2808 -264 2844 -252
rect 2856 -264 2868 -252
rect 2880 -264 2916 -252
rect 2928 -264 2940 -252
rect 2952 -264 2988 -252
rect -1020 -288 2988 -264
rect -1020 -300 -996 -288
rect -984 -300 -972 -288
rect -960 -300 -948 -288
rect -936 -300 -924 -288
rect -912 -300 -900 -288
rect -888 -300 -876 -288
rect -864 -300 -852 -288
rect -840 -300 -828 -288
rect -816 -300 -804 -288
rect -792 -300 -780 -288
rect -768 -300 -756 -288
rect -744 -300 -732 -288
rect -720 -300 -708 -288
rect -696 -300 -684 -288
rect -672 -300 -660 -288
rect -648 -300 -636 -288
rect -624 -300 -612 -288
rect -600 -300 -588 -288
rect -576 -300 -564 -288
rect -552 -300 -540 -288
rect -528 -300 -516 -288
rect -504 -300 -492 -288
rect -480 -300 -468 -288
rect -456 -300 -444 -288
rect -432 -300 -420 -288
rect -408 -300 -396 -288
rect -384 -300 -372 -288
rect -360 -300 -348 -288
rect -336 -300 -324 -288
rect -312 -300 -300 -288
rect -288 -300 -276 -288
rect -264 -300 -252 -288
rect -240 -300 -228 -288
rect -216 -300 -204 -288
rect -192 -300 -180 -288
rect -168 -300 -156 -288
rect -144 -300 -132 -288
rect -120 -300 -108 -288
rect -96 -300 -84 -288
rect -72 -300 -60 -288
rect -48 -300 -36 -288
rect -24 -300 -12 -288
rect 0 -300 12 -288
rect 24 -300 36 -288
rect 48 -300 60 -288
rect 72 -300 84 -288
rect 96 -300 108 -288
rect 120 -300 132 -288
rect 144 -300 156 -288
rect 168 -300 180 -288
rect 192 -300 204 -288
rect 216 -300 228 -288
rect 240 -300 252 -288
rect 264 -300 276 -288
rect 288 -300 300 -288
rect 312 -300 324 -288
rect 336 -300 348 -288
rect 360 -300 372 -288
rect 384 -300 396 -288
rect 408 -300 420 -288
rect 432 -300 444 -288
rect 456 -300 468 -288
rect 480 -300 492 -288
rect 504 -300 516 -288
rect 528 -300 540 -288
rect 552 -300 564 -288
rect 576 -300 588 -288
rect 600 -300 612 -288
rect 624 -300 636 -288
rect 648 -300 660 -288
rect 672 -300 684 -288
rect 696 -300 708 -288
rect 720 -300 732 -288
rect 744 -300 756 -288
rect 768 -300 780 -288
rect 792 -300 804 -288
rect 816 -300 828 -288
rect 840 -300 852 -288
rect 864 -300 876 -288
rect 888 -300 900 -288
rect 912 -300 924 -288
rect 936 -300 948 -288
rect 960 -300 972 -288
rect 984 -300 996 -288
rect 1008 -300 1020 -288
rect 1032 -300 1044 -288
rect 1056 -300 1068 -288
rect 1080 -300 1092 -288
rect 1104 -300 1116 -288
rect 1128 -300 1140 -288
rect 1152 -300 1164 -288
rect 1176 -300 1188 -288
rect 1200 -300 1212 -288
rect 1224 -300 1236 -288
rect 1248 -300 1260 -288
rect 1272 -300 1284 -288
rect 1296 -300 1308 -288
rect 1320 -300 1332 -288
rect 1344 -300 1356 -288
rect 1368 -300 1380 -288
rect 1392 -300 1404 -288
rect 1416 -300 1428 -288
rect 1440 -300 1452 -288
rect 1464 -300 1476 -288
rect 1488 -300 1500 -288
rect 1512 -300 1524 -288
rect 1536 -300 1548 -288
rect 1560 -300 1572 -288
rect 1584 -300 1596 -288
rect 1608 -300 1620 -288
rect 1632 -300 1644 -288
rect 1656 -300 1668 -288
rect 1680 -300 1692 -288
rect 1704 -300 1716 -288
rect 1728 -300 1740 -288
rect 1752 -300 1764 -288
rect 1776 -300 1788 -288
rect 1800 -300 1812 -288
rect 1824 -300 1836 -288
rect 1848 -300 1860 -288
rect 1872 -300 1884 -288
rect 1896 -300 1908 -288
rect 1920 -300 1932 -288
rect 1944 -300 1956 -288
rect 1968 -300 1980 -288
rect 1992 -300 2004 -288
rect 2016 -300 2028 -288
rect 2040 -300 2052 -288
rect 2064 -300 2076 -288
rect 2088 -300 2100 -288
rect 2112 -300 2124 -288
rect 2136 -300 2148 -288
rect 2160 -300 2172 -288
rect 2184 -300 2196 -288
rect 2208 -300 2220 -288
rect 2232 -300 2244 -288
rect 2256 -300 2268 -288
rect 2280 -300 2292 -288
rect 2304 -300 2316 -288
rect 2328 -300 2340 -288
rect 2352 -300 2364 -288
rect 2376 -300 2388 -288
rect 2400 -300 2412 -288
rect 2424 -300 2436 -288
rect 2448 -300 2460 -288
rect 2472 -300 2484 -288
rect 2496 -300 2508 -288
rect 2520 -300 2532 -288
rect 2544 -300 2556 -288
rect 2568 -300 2580 -288
rect 2592 -300 2604 -288
rect 2616 -300 2628 -288
rect 2640 -300 2652 -288
rect 2664 -300 2676 -288
rect 2688 -300 2700 -288
rect 2712 -300 2724 -288
rect 2736 -300 2748 -288
rect 2760 -300 2772 -288
rect 2784 -300 2796 -288
rect 2808 -300 2820 -288
rect 2832 -300 2844 -288
rect 2856 -300 2868 -288
rect 2880 -300 2892 -288
rect 2904 -300 2916 -288
rect 2928 -300 2940 -288
rect 2952 -300 2988 -288
rect -1020 -324 2988 -300
rect -1020 -336 -996 -324
rect -984 -336 -972 -324
rect -960 -336 -948 -324
rect -936 -336 -924 -324
rect -912 -336 -900 -324
rect -888 -336 -876 -324
rect -864 -336 -852 -324
rect -840 -336 -828 -324
rect -816 -336 -804 -324
rect -792 -336 -780 -324
rect -768 -336 -756 -324
rect -744 -336 -732 -324
rect -720 -336 -708 -324
rect -696 -336 -684 -324
rect -672 -336 -660 -324
rect -648 -336 -636 -324
rect -624 -336 -612 -324
rect -600 -336 -588 -324
rect -576 -336 -564 -324
rect -552 -336 -540 -324
rect -528 -336 -516 -324
rect -504 -336 -492 -324
rect -480 -336 -468 -324
rect -456 -336 -444 -324
rect -432 -336 -420 -324
rect -408 -336 -396 -324
rect -384 -336 -372 -324
rect -360 -336 -348 -324
rect -336 -336 -324 -324
rect -312 -336 -300 -324
rect -288 -336 -276 -324
rect -264 -336 -252 -324
rect -240 -336 -228 -324
rect -216 -336 -204 -324
rect -192 -336 -180 -324
rect -168 -336 -156 -324
rect -144 -336 -132 -324
rect -120 -336 -108 -324
rect -96 -336 -84 -324
rect -72 -336 -60 -324
rect -48 -336 -36 -324
rect -24 -336 -12 -324
rect 0 -336 12 -324
rect 24 -336 36 -324
rect 48 -336 60 -324
rect 72 -336 84 -324
rect 96 -336 108 -324
rect 120 -336 132 -324
rect 144 -336 156 -324
rect 168 -336 180 -324
rect 192 -336 204 -324
rect 216 -336 228 -324
rect 240 -336 252 -324
rect 264 -336 276 -324
rect 288 -336 300 -324
rect 312 -336 324 -324
rect 336 -336 348 -324
rect 360 -336 372 -324
rect 384 -336 396 -324
rect 408 -336 420 -324
rect 432 -336 444 -324
rect 456 -336 468 -324
rect 480 -336 492 -324
rect 504 -336 516 -324
rect 528 -336 540 -324
rect 552 -336 564 -324
rect 576 -336 588 -324
rect 600 -336 612 -324
rect 624 -336 636 -324
rect 648 -336 660 -324
rect 672 -336 684 -324
rect 696 -336 708 -324
rect 720 -336 732 -324
rect 744 -336 756 -324
rect 768 -336 780 -324
rect 792 -336 804 -324
rect 816 -336 828 -324
rect 840 -336 852 -324
rect 864 -336 876 -324
rect 888 -336 900 -324
rect 912 -336 924 -324
rect 936 -336 948 -324
rect 960 -336 972 -324
rect 984 -336 996 -324
rect 1008 -336 1020 -324
rect 1032 -336 1044 -324
rect 1056 -336 1068 -324
rect 1080 -336 1092 -324
rect 1104 -336 1116 -324
rect 1128 -336 1140 -324
rect 1152 -336 1164 -324
rect 1176 -336 1188 -324
rect 1200 -336 1212 -324
rect 1224 -336 1236 -324
rect 1248 -336 1260 -324
rect 1272 -336 1284 -324
rect 1296 -336 1308 -324
rect 1320 -336 1332 -324
rect 1344 -336 1356 -324
rect 1368 -336 1380 -324
rect 1392 -336 1404 -324
rect 1416 -336 1428 -324
rect 1440 -336 1452 -324
rect 1464 -336 1476 -324
rect 1488 -336 1500 -324
rect 1512 -336 1524 -324
rect 1536 -336 1548 -324
rect 1560 -336 1572 -324
rect 1584 -336 1596 -324
rect 1608 -336 1620 -324
rect 1632 -336 1644 -324
rect 1656 -336 1668 -324
rect 1680 -336 1692 -324
rect 1704 -336 1716 -324
rect 1728 -336 1740 -324
rect 1752 -336 1764 -324
rect 1776 -336 1788 -324
rect 1800 -336 1812 -324
rect 1824 -336 1836 -324
rect 1848 -336 1860 -324
rect 1872 -336 1884 -324
rect 1896 -336 1908 -324
rect 1920 -336 1932 -324
rect 1944 -336 1956 -324
rect 1968 -336 1980 -324
rect 1992 -336 2004 -324
rect 2016 -336 2028 -324
rect 2040 -336 2052 -324
rect 2064 -336 2076 -324
rect 2088 -336 2100 -324
rect 2112 -336 2124 -324
rect 2136 -336 2148 -324
rect 2160 -336 2172 -324
rect 2184 -336 2196 -324
rect 2208 -336 2220 -324
rect 2232 -336 2244 -324
rect 2256 -336 2268 -324
rect 2280 -336 2292 -324
rect 2304 -336 2316 -324
rect 2328 -336 2340 -324
rect 2352 -336 2364 -324
rect 2376 -336 2388 -324
rect 2400 -336 2412 -324
rect 2424 -336 2436 -324
rect 2448 -336 2460 -324
rect 2472 -336 2484 -324
rect 2496 -336 2508 -324
rect 2520 -336 2532 -324
rect 2544 -336 2556 -324
rect 2568 -336 2580 -324
rect 2592 -336 2604 -324
rect 2616 -336 2628 -324
rect 2640 -336 2652 -324
rect 2664 -336 2676 -324
rect 2688 -336 2700 -324
rect 2712 -336 2724 -324
rect 2736 -336 2748 -324
rect 2760 -336 2772 -324
rect 2784 -336 2796 -324
rect 2808 -336 2820 -324
rect 2832 -336 2844 -324
rect 2856 -336 2868 -324
rect 2880 -336 2892 -324
rect 2904 -336 2916 -324
rect 2928 -336 2940 -324
rect 2952 -336 2988 -324
rect -1020 -360 2988 -336
rect -1020 -372 -996 -360
rect -984 -372 -972 -360
rect -960 -372 -948 -360
rect -936 -372 -924 -360
rect -912 -372 -900 -360
rect -888 -372 -876 -360
rect -864 -372 -852 -360
rect -840 -372 -828 -360
rect -816 -372 -804 -360
rect -792 -372 -780 -360
rect -768 -372 -756 -360
rect -744 -372 -732 -360
rect -720 -372 -708 -360
rect -696 -372 -684 -360
rect -672 -372 -660 -360
rect -648 -372 -636 -360
rect -624 -372 -612 -360
rect -600 -372 -588 -360
rect -576 -372 -564 -360
rect -552 -372 -540 -360
rect -528 -372 -516 -360
rect -504 -372 -492 -360
rect -480 -372 -468 -360
rect -456 -372 -444 -360
rect -432 -372 -420 -360
rect -408 -372 -396 -360
rect -384 -372 -372 -360
rect -360 -372 -348 -360
rect -336 -372 -324 -360
rect -312 -372 -300 -360
rect -288 -372 -276 -360
rect -264 -372 -252 -360
rect -240 -372 -228 -360
rect -216 -372 -204 -360
rect -192 -372 -180 -360
rect -168 -372 -156 -360
rect -144 -372 -132 -360
rect -120 -372 -108 -360
rect -96 -372 -84 -360
rect -72 -372 -60 -360
rect -48 -372 -36 -360
rect -24 -372 -12 -360
rect 0 -372 12 -360
rect 24 -372 36 -360
rect 48 -372 60 -360
rect 72 -372 84 -360
rect 96 -372 108 -360
rect 120 -372 132 -360
rect 144 -372 156 -360
rect 168 -372 180 -360
rect 192 -372 204 -360
rect 216 -372 228 -360
rect 240 -372 252 -360
rect 264 -372 276 -360
rect 288 -372 300 -360
rect 312 -372 324 -360
rect 336 -372 348 -360
rect 360 -372 372 -360
rect 384 -372 396 -360
rect 408 -372 420 -360
rect 432 -372 444 -360
rect 456 -372 468 -360
rect 480 -372 492 -360
rect 504 -372 516 -360
rect 528 -372 540 -360
rect 552 -372 564 -360
rect 576 -372 588 -360
rect 600 -372 612 -360
rect 624 -372 636 -360
rect 648 -372 660 -360
rect 672 -372 684 -360
rect 696 -372 708 -360
rect 720 -372 732 -360
rect 744 -372 756 -360
rect 768 -372 780 -360
rect 792 -372 804 -360
rect 816 -372 828 -360
rect 840 -372 852 -360
rect 864 -372 876 -360
rect 888 -372 900 -360
rect 912 -372 924 -360
rect 936 -372 948 -360
rect 960 -372 972 -360
rect 984 -372 996 -360
rect 1008 -372 1020 -360
rect 1032 -372 1044 -360
rect 1056 -372 1068 -360
rect 1080 -372 1092 -360
rect 1104 -372 1116 -360
rect 1128 -372 1140 -360
rect 1152 -372 1164 -360
rect 1176 -372 1188 -360
rect 1200 -372 1212 -360
rect 1224 -372 1236 -360
rect 1248 -372 1260 -360
rect 1272 -372 1284 -360
rect 1296 -372 1308 -360
rect 1320 -372 1332 -360
rect 1344 -372 1356 -360
rect 1368 -372 1380 -360
rect 1392 -372 1404 -360
rect 1416 -372 1428 -360
rect 1440 -372 1452 -360
rect 1464 -372 1476 -360
rect 1488 -372 1500 -360
rect 1512 -372 1524 -360
rect 1536 -372 1548 -360
rect 1560 -372 1572 -360
rect 1584 -372 1596 -360
rect 1608 -372 1620 -360
rect 1632 -372 1644 -360
rect 1656 -372 1668 -360
rect 1680 -372 1692 -360
rect 1704 -372 1716 -360
rect 1728 -372 1740 -360
rect 1752 -372 1764 -360
rect 1776 -372 1788 -360
rect 1800 -372 1812 -360
rect 1824 -372 1836 -360
rect 1848 -372 1860 -360
rect 1872 -372 1884 -360
rect 1896 -372 1908 -360
rect 1920 -372 1932 -360
rect 1944 -372 1956 -360
rect 1968 -372 1980 -360
rect 1992 -372 2004 -360
rect 2016 -372 2028 -360
rect 2040 -372 2052 -360
rect 2064 -372 2076 -360
rect 2088 -372 2100 -360
rect 2112 -372 2124 -360
rect 2136 -372 2148 -360
rect 2160 -372 2172 -360
rect 2184 -372 2196 -360
rect 2208 -372 2220 -360
rect 2232 -372 2244 -360
rect 2256 -372 2268 -360
rect 2280 -372 2292 -360
rect 2304 -372 2316 -360
rect 2328 -372 2340 -360
rect 2352 -372 2364 -360
rect 2376 -372 2388 -360
rect 2400 -372 2412 -360
rect 2424 -372 2436 -360
rect 2448 -372 2460 -360
rect 2472 -372 2484 -360
rect 2496 -372 2508 -360
rect 2520 -372 2532 -360
rect 2544 -372 2556 -360
rect 2568 -372 2580 -360
rect 2592 -372 2604 -360
rect 2616 -372 2628 -360
rect 2640 -372 2652 -360
rect 2664 -372 2676 -360
rect 2688 -372 2700 -360
rect 2712 -372 2724 -360
rect 2736 -372 2748 -360
rect 2760 -372 2772 -360
rect 2784 -372 2796 -360
rect 2808 -372 2820 -360
rect 2832 -372 2844 -360
rect 2856 -372 2868 -360
rect 2880 -372 2892 -360
rect 2904 -372 2916 -360
rect 2928 -372 2940 -360
rect 2952 -372 2988 -360
rect -1020 -396 2988 -372
use manfvieru_cell  manfvieru_cell_0
timestamp 1664997892
transform 1 0 252 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_1
timestamp 1664997892
transform 1 0 372 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_2
timestamp 1664997892
transform 1 0 492 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_3
timestamp 1664997892
transform 1 0 612 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_4
timestamp 1664997892
transform 1 0 732 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_5
timestamp 1664997892
transform 1 0 852 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_6
timestamp 1664997892
transform 1 0 972 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_7
timestamp 1664997892
transform 1 0 1092 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_8
timestamp 1664997892
transform 1 0 1212 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_9
timestamp 1664997892
transform 1 0 1332 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_10
timestamp 1664997892
transform 1 0 1452 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_11
timestamp 1664997892
transform -1 0 264 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_12
timestamp 1664997892
transform -1 0 384 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_13
timestamp 1664997892
transform -1 0 -1176 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_14
timestamp 1664997892
transform 1 0 -228 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_15
timestamp 1664997892
transform -1 0 -1296 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_16
timestamp 1664997892
transform 1 0 -108 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_17
timestamp 1664997892
transform -1 0 2424 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_18
timestamp 1664997892
transform 1 0 3492 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_19
timestamp 1664997892
transform -1 0 2304 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_20
timestamp 1664997892
transform -1 0 1944 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_21
timestamp 1664997892
transform 1 0 3372 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_22
timestamp 1664997892
transform -1 0 1704 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_23
timestamp 1664997892
transform -1 0 1824 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_24
timestamp 1664997892
transform -1 0 1464 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_25
timestamp 1664997892
transform -1 0 1584 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_26
timestamp 1664997892
transform -1 0 1224 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_27
timestamp 1664997892
transform -1 0 1344 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_28
timestamp 1664997892
transform -1 0 1104 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_29
timestamp 1664997892
transform -1 0 984 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_30
timestamp 1664997892
transform -1 0 744 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_31
timestamp 1664997892
transform -1 0 864 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_32
timestamp 1664997892
transform 1 0 1812 0 1 -36
box -720 -132 -588 708
use manfvieru_cell  manfvieru_cell_33
timestamp 1664997892
transform 1 0 1932 0 1 -36
box -720 -132 -588 708
use manfvieru_edge  manfvieru_edge_0
timestamp 1664998004
transform 1 0 -276 0 1 -36
box -756 -132 -660 708
use manfvieru_edge  manfvieru_edge_1
timestamp 1664998004
transform -1 0 2472 0 1 -36
box -756 -132 -660 708
<< labels >>
rlabel metal3 -1044 -168 -1032 -108 0 gnd
port 9 nsew
rlabel metal3 -1044 -48 -1032 -36 0 om
port 4 nsew
rlabel metal3 -1044 -12 -1032 0 0 xp
rlabel metal3 -1044 588 -1032 648 0 vdd
port 5 nsew
rlabel metal3 -1044 516 -1032 528 0 gp
port 6 nsew
rlabel metal3 -1044 384 -1032 396 0 bp
port 7 nsew
rlabel metal3 -1044 540 -1032 552 0 vreg
port 8 nsew
rlabel metal3 -1044 216 -1032 228 0 im
port 2 nsew
rlabel metal3 -1044 336 -1032 348 0 op
port 3 nsew
rlabel metal3 -1044 300 -1032 312 0 xm
rlabel metal3 -1044 168 -1032 180 0 x
rlabel metal3 -1044 72 -1032 84 0 ip
port 1 nsew
rlabel metal3 -1044 120 -1032 132 0 y
<< end >>
