.subckt pch6 d g s b
x0 d g s b pmos_6p0 w=1.8u l=0.6u
x1 d g s b pmos_6p0 w=1.8u l=0.6u
.ends

.subckt nch6 d g s b
x0 x g s b nmos_6p0 w=1.8u l=0.6u
x1 d g x b nmos_6p0 w=1.8u l=0.6u
.ends

.subckt pch3 d g s b
x0 d g s b pmos_3p3 w=1.5u l=0.6u
x1 d g s b pmos_3p3 w=1.5u l=0.6u
.ends

.subckt nch3 d g s b
x0 x g s b nmos_3p3 w=1.8u l=0.6u
x1 d g x b nmos_3p3 w=1.8u l=0.6u
.ends

.subckt inv0 in out vdd gp bp vreg gnd
XV  vreg gp vdd  vdd pch6
XP  out  in vreg bp  pch3
XN  out  in gnd  gnd nch3
.ends

.subckt qref p ref m lo
XPV1 x   x   p   p   pmos_6p0 w=6.0u l=6.0u
XPV2 ref ref x   x   pmos_6p0 w=6.0u l=6.0u
XPV3 y   y   ref ref pmos_6p0 w=6.0u l=6.0u
XPV4 m   lo  y   y   pmos_6p0 w=6.0u l=6.0u
.ends

.subckt inv_bias ib vdd gp bp vreg gnd
XP1a vreg gp  vdd  vdd pch6
XP1b q    q   vreg bp  pch3
XN1c q    q   gnd  gnd nch3

XP2a z    z    vdd  vdd pch6
XN2b z    vreg y    gnd nch6
XN2c y    q    gnd  gnd nch3

XP3a gp   z    vdd  vdd pch6
XN3b gp   vreg x    gnd nch6
XN3c x    ib   gnd  gnd nch6

XNV4 ib   ib  gnd  gnd nch6

xref vreg ref gnd  gnd qref

XP5a vreg gp  vdd  vdd pch6
XP5b bp0  ref vreg bp  pch3
XN5c bp0  ref gnd  gnd nch3

XP6a bp   gp0 vdd  vdd pch6
XP6b gnd  bp0 bp   bp  pch3
XN6c gnd  bp0 gnd  gnd nch3

XPV7 gp0  gp0 vdd  vdd pch6
XNV7 gp0  ib  gnd  gnd nch6


cc vdd gp 10f

.ends
