* NGSPICE file created from nautavieru.ext - technology: gf180mcuC

.subckt nautavieru_cell inl inr out gp vreg op xm im ip xp om x vdd gnd bp
X0 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X1 vreg inr out bp pmos_3p3 w=1.5u l=0.6u
X2 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X3 dr inr out gnd nmos_3p3 w=1.8u l=0.6u
X4 dl inl gnd gnd nmos_3p3 w=1.8u l=0.6u
X5 out inr vreg bp pmos_3p3 w=1.5u l=0.6u
X6 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X7 vreg inl out bp pmos_3p3 w=1.5u l=0.6u
X8 gnd inr dr gnd nmos_3p3 w=1.8u l=0.6u
X9 out inl dl gnd nmos_3p3 w=1.8u l=0.6u
X10 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X11 out inl vreg bp pmos_3p3 w=1.5u l=0.6u
C0 out vreg 0.78fF
C1 inl om 0.18fF
C2 op inl 0.20fF
C3 vdd vreg 1.41fF
C4 out bp 0.15fF
C5 bp vreg 0.92fF
C6 inr om 0.18fF
C7 op inr 0.20fF
C8 inl inr 0.60fF
C9 xp om 1.35fF
C10 out om 0.12fF
C11 op out 0.12fF
C12 inl out 0.17fF
C13 gp vreg 1.98fF
C14 vdd gp 0.66fF
C15 inl bp 0.32fF
C16 inr out 0.20fF
C17 xm op 1.35fF
C18 inr bp 0.32fF
C19 out gnd 1.64fF
C20 inr gnd 2.31fF
C21 inl gnd 2.32fF
C22 vreg gnd 0.72fF
C23 gp gnd 1.56fF
C24 bp gnd 6.58fF
C25 vdd gnd 6.08fF
C26 dr gnd 0.18fF
C27 dl gnd 0.18fF
.ends

.subckt nautavieru_edge gp vreg im ip xm op xp om x vdd gnd bp
X0 gnd lo lo gnd nmos_3p3 w=1.8u l=0.6u
X1 vdd hih hih vdd pmos_6p0 w=1.8u l=0.6u
X2 vreg hi hi bp pmos_3p3 w=1.5u l=0.6u
C0 hi vreg 0.11fF
C1 gp vreg 1.01fF
C2 bp vreg 0.23fF
C3 hi bp 0.28fF
C4 op xm 0.98fF
C5 om xp 0.98fF
C6 hih vdd 0.45fF
C7 vdd vreg 0.22fF
C8 vreg gnd 0.44fF
C9 bp gnd 4.35fF
C10 vdd gnd 4.01fF
C11 lo gnd 0.84fF
C12 hi gnd 0.46fF
C13 hih gnd 0.46fF
.ends

.subckt nautavieru ip im op om vdd gp bp vreg gnd
Xnautavieru_cell_16 ip xm xm gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_26 x x xm gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_27 ip ip om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_15 ip ip om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_17 ip xp xm gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_28 xp xp om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_18 xm im xp gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_29 im im op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_19 xp im xp gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_edge_0 gp vreg im ip xm op xp om x vdd gnd bp nautavieru_edge
Xnautavieru_edge_1 gp vreg im ip xm op xp om x vdd gnd bp nautavieru_edge
Xnautavieru_cell_0 ip xm xm gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_1 xm im xp gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_2 ip xp xm gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_3 xp im xp gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_4 xp xp om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_5 xm xm op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_7 x op x gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_6 om x x gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_8 x x xp gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_9 xm xm op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_30 im im op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_20 xp xp om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_31 ip ip om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_21 xm xm op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_10 xp xp om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_22 om x x gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_11 x x xm gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_23 x x xp gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_12 ip ip om gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_24 x op x gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_13 im im op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_25 xm xm op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
Xnautavieru_cell_14 im im op gp vreg op xm im ip xp om x vdd gnd bp nautavieru_cell
X0 om xp mim_2p0fF c_width=199.2u c_length=7.2u
X1 op xm mim_2p0fF c_width=199.2u c_length=7.2u
C0 xp vreg 0.19fF
C1 op im 0.61fF
C2 im x 0.18fF
C3 op ip 0.73fF
C4 xm im 0.13fF
C5 x ip 0.20fF
C6 op om 0.48fF
C7 im xp 1.91fF
C8 xm ip 0.99fF
C9 x om 0.68fF
C10 ip xp 1.18fF
C11 xm om 1.64fF
C12 xp om 47.50fF
C13 gp vdd 0.30fF
C14 op vdd 4.12fF
C15 gp op 0.63fF
C16 xm vdd 5.00fF
C17 gp xm 0.59fF
C18 om vreg 0.16fF
C19 op x 1.37fF
C20 xm op 47.73fF
C21 op bp 0.13fF
C22 op xp 0.76fF
C23 im ip 1.82fF
C24 xm x 1.23fF
C25 x xp 0.53fF
C26 im om 0.87fF
C27 xm xp 3.05fF
C28 vreg vdd 0.75fF
C29 ip om 0.94fF
C30 gp vreg -2.33fF
C31 op vreg 1.04fF
C32 x vreg 0.16fF
C33 xm vreg 1.06fF
C34 vreg bp 0.11fF
C35 bp gnd 195.36fF
C36 vdd gnd 173.19fF
C37 om gnd 68.09fF
C38 xp gnd 47.10fF
C39 ip gnd 50.03fF
C40 x gnd 56.38fF
C41 im gnd 48.37fF
C42 op gnd 53.53fF
C43 xm gnd 42.27fF
C44 gp gnd 44.32fF
C45 vreg gnd 8.33fF
.ends

