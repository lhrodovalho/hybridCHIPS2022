* NGSPICE file created from manfvieru.ext - technology: gf180mcuC

.subckt manfvieru_edge gp vreg im ip xm op xp om x y vdd gnd bp
X0 vreg hi hi bp pmos_3p3 w=1.5u l=0.6u
X1 gnd lo lo gnd nmos_3p3 w=1.8u l=0.6u
X2 vdd hih hih vdd pmos_6p0 w=1.8u l=0.6u
C0 vreg gp 1.01fF
C1 xm op 0.98fF
C2 vdd hih 0.45fF
C3 om xp 0.98fF
C4 vreg bp 0.23fF
C5 hi bp 0.28fF
C6 vreg vdd 0.22fF
C7 vreg hi 0.11fF
C8 vreg gnd 0.44fF
C9 bp gnd 4.35fF
C10 vdd gnd 4.01fF
C11 lo gnd 0.84fF
C12 hi gnd 0.46fF
C13 hih gnd 0.46fF
.ends

.subckt manfvieru_cell inl inr out gp vreg op xm im ip xp om x y vdd gnd bp
X0 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X1 out inl vreg bp pmos_3p3 w=1.5u l=0.6u
X2 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X3 vdd gp vreg vdd pmos_6p0 w=1.8u l=0.6u
X4 dr inr out gnd nmos_3p3 w=1.8u l=0.6u
X5 dl inl gnd gnd nmos_3p3 w=1.8u l=0.6u
X6 vreg inr out bp pmos_3p3 w=1.5u l=0.6u
X7 gnd inr dr gnd nmos_3p3 w=1.8u l=0.6u
X8 out inl dl gnd nmos_3p3 w=1.8u l=0.6u
X9 vreg gp vdd vdd pmos_6p0 w=1.8u l=0.6u
X10 out inr vreg bp pmos_3p3 w=1.5u l=0.6u
X11 vreg inl out bp pmos_3p3 w=1.5u l=0.6u
C0 op xm 1.35fF
C1 bp out 0.15fF
C2 op out 0.12fF
C3 om out 0.12fF
C4 inl bp 0.32fF
C5 inl op 0.20fF
C6 om inl 0.18fF
C7 out inr 0.20fF
C8 inl inr 0.64fF
C9 vreg vdd 1.41fF
C10 vdd gp 0.66fF
C11 om xp 1.35fF
C12 vreg gp 1.98fF
C13 vreg out 0.78fF
C14 bp inr 0.32fF
C15 op inr 0.20fF
C16 om inr 0.18fF
C17 inl out 0.18fF
C18 vreg bp 0.92fF
C19 out gnd 1.80fF
C20 inr gnd 2.38fF
C21 inl gnd 2.39fF
C22 vreg gnd 0.72fF
C23 gp gnd 1.56fF
C24 bp gnd 6.58fF
C25 vdd gnd 6.08fF
C26 dr gnd 0.18fF
C27 dl gnd 0.18fF
.ends

.subckt manfvieru ip im op om vdd gp bp vreg gnd
Xmanfvieru_edge_0 gp vreg im ip xm op xp om x y vdd gnd bp manfvieru_edge
Xmanfvieru_edge_1 gp vreg im ip xm op xp om x y vdd gnd bp manfvieru_edge
Xmanfvieru_cell_0 im y xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_1 y ip xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_2 xp x x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_30 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_3 x om y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_20 im y xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_31 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_4 y y y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_21 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_32 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_10 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_5 op x y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_22 xp x x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_33 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_11 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_7 ip y xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_6 x xm x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_23 y ip xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_12 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_8 y im xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_24 y y y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_9 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_13 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_25 x om y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_14 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_27 op x y gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_26 x xm x gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_15 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_16 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_17 xp ip om gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_28 ip y xm gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_18 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_29 y im xp gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
Xmanfvieru_cell_19 im xm op gp vreg op xm im ip xp om x y vdd gnd bp manfvieru_cell
X0 om xp mim_2p0fF c_width=199.2u c_length=7.2u
X1 op xm mim_2p0fF c_width=199.2u c_length=7.2u
C0 vreg x 0.13fF
C1 xm op 52.52fF
C2 om op 0.43fF
C3 xm x 0.20fF
C4 op im 0.52fF
C5 xp bp 0.11fF
C6 vreg vdd 0.78fF
C7 om x 0.41fF
C8 im x 0.15fF
C9 xm ip 1.12fF
C10 op y 1.33fF
C11 om ip 0.66fF
C12 x y 0.53fF
C13 op xp 0.67fF
C14 im ip 3.37fF
C15 xm vdd 5.43fF
C16 x xp 0.29fF
C17 y ip 0.20fF
C18 vreg xm 1.31fF
C19 gp op 0.65fF
C20 ip xp 1.04fF
C21 om vreg 0.16fF
C22 op bp 0.13fF
C23 vreg y 0.20fF
C24 om xm 0.66fF
C25 xm im 0.11fF
C26 vreg xp 0.14fF
C27 gp vdd 0.27fF
C28 om im 1.05fF
C29 op x 0.28fF
C30 xm y 0.36fF
C31 gp vreg -2.47fF
C32 om y 1.64fF
C33 im y 0.15fF
C34 xm xp 0.52fF
C35 op ip 0.71fF
C36 om xp 52.23fF
C37 x ip 0.37fF
C38 im xp 2.13fF
C39 gp xm 0.72fF
C40 op vdd 4.12fF
C41 y xp 0.72fF
C42 vreg op 1.05fF
C43 bp gnd 207.63fF
C44 vdd gnd 183.59fF
C45 om gnd 71.62fF
C46 xp gnd 41.51fF
C47 ip gnd 52.08fF
C48 y gnd 63.08fF
C49 x gnd 49.40fF
C50 im gnd 52.06fF
C51 op gnd 56.87fF
C52 xm gnd 35.93fF
C53 vreg gnd 9.16fF
C54 gp gnd 47.13fF
.ends

